magic
tech sky130A
magscale 1 2
timestamp 1754688798
<< error_p >>
rect -29 210 29 216
rect -29 176 -17 210
rect -29 170 29 176
<< nwell >>
rect -109 -263 109 229
<< pmos >>
rect -15 -201 15 129
<< pdiff >>
rect -73 117 -15 129
rect -73 -189 -61 117
rect -27 -189 -15 117
rect -73 -201 -15 -189
rect 15 117 73 129
rect 15 -189 27 117
rect 61 -189 73 117
rect 15 -201 73 -189
<< pdiffc >>
rect -61 -189 -27 117
rect 27 -189 61 117
<< poly >>
rect -33 210 33 226
rect -33 176 -17 210
rect 17 176 33 210
rect -33 160 33 176
rect -15 129 15 160
rect -15 -227 15 -201
<< polycont >>
rect -17 176 17 210
<< locali >>
rect -33 176 -17 210
rect 17 176 33 210
rect -61 117 -27 133
rect -61 -205 -27 -189
rect 27 117 61 133
rect 27 -205 61 -189
<< viali >>
rect -17 176 17 210
rect -61 -189 -27 117
rect 27 -189 61 117
<< metal1 >>
rect -29 210 29 216
rect -29 176 -17 210
rect 17 176 29 210
rect -29 170 29 176
rect -67 117 -21 129
rect -67 -189 -61 117
rect -27 -189 -21 117
rect -67 -201 -21 -189
rect 21 117 67 129
rect 21 -189 27 117
rect 61 -189 67 117
rect 21 -201 67 -189
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.65 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1754900058
<< metal3 >>
rect -686 84332 686 84360
rect -686 83308 602 84332
rect 666 83308 686 84332
rect -686 83280 686 83308
rect -686 83012 686 83040
rect -686 81988 602 83012
rect 666 81988 686 83012
rect -686 81960 686 81988
rect -686 81692 686 81720
rect -686 80668 602 81692
rect 666 80668 686 81692
rect -686 80640 686 80668
rect -686 80372 686 80400
rect -686 79348 602 80372
rect 666 79348 686 80372
rect -686 79320 686 79348
rect -686 79052 686 79080
rect -686 78028 602 79052
rect 666 78028 686 79052
rect -686 78000 686 78028
rect -686 77732 686 77760
rect -686 76708 602 77732
rect 666 76708 686 77732
rect -686 76680 686 76708
rect -686 76412 686 76440
rect -686 75388 602 76412
rect 666 75388 686 76412
rect -686 75360 686 75388
rect -686 75092 686 75120
rect -686 74068 602 75092
rect 666 74068 686 75092
rect -686 74040 686 74068
rect -686 73772 686 73800
rect -686 72748 602 73772
rect 666 72748 686 73772
rect -686 72720 686 72748
rect -686 72452 686 72480
rect -686 71428 602 72452
rect 666 71428 686 72452
rect -686 71400 686 71428
rect -686 71132 686 71160
rect -686 70108 602 71132
rect 666 70108 686 71132
rect -686 70080 686 70108
rect -686 69812 686 69840
rect -686 68788 602 69812
rect 666 68788 686 69812
rect -686 68760 686 68788
rect -686 68492 686 68520
rect -686 67468 602 68492
rect 666 67468 686 68492
rect -686 67440 686 67468
rect -686 67172 686 67200
rect -686 66148 602 67172
rect 666 66148 686 67172
rect -686 66120 686 66148
rect -686 65852 686 65880
rect -686 64828 602 65852
rect 666 64828 686 65852
rect -686 64800 686 64828
rect -686 64532 686 64560
rect -686 63508 602 64532
rect 666 63508 686 64532
rect -686 63480 686 63508
rect -686 63212 686 63240
rect -686 62188 602 63212
rect 666 62188 686 63212
rect -686 62160 686 62188
rect -686 61892 686 61920
rect -686 60868 602 61892
rect 666 60868 686 61892
rect -686 60840 686 60868
rect -686 60572 686 60600
rect -686 59548 602 60572
rect 666 59548 686 60572
rect -686 59520 686 59548
rect -686 59252 686 59280
rect -686 58228 602 59252
rect 666 58228 686 59252
rect -686 58200 686 58228
rect -686 57932 686 57960
rect -686 56908 602 57932
rect 666 56908 686 57932
rect -686 56880 686 56908
rect -686 56612 686 56640
rect -686 55588 602 56612
rect 666 55588 686 56612
rect -686 55560 686 55588
rect -686 55292 686 55320
rect -686 54268 602 55292
rect 666 54268 686 55292
rect -686 54240 686 54268
rect -686 53972 686 54000
rect -686 52948 602 53972
rect 666 52948 686 53972
rect -686 52920 686 52948
rect -686 52652 686 52680
rect -686 51628 602 52652
rect 666 51628 686 52652
rect -686 51600 686 51628
rect -686 51332 686 51360
rect -686 50308 602 51332
rect 666 50308 686 51332
rect -686 50280 686 50308
rect -686 50012 686 50040
rect -686 48988 602 50012
rect 666 48988 686 50012
rect -686 48960 686 48988
rect -686 48692 686 48720
rect -686 47668 602 48692
rect 666 47668 686 48692
rect -686 47640 686 47668
rect -686 47372 686 47400
rect -686 46348 602 47372
rect 666 46348 686 47372
rect -686 46320 686 46348
rect -686 46052 686 46080
rect -686 45028 602 46052
rect 666 45028 686 46052
rect -686 45000 686 45028
rect -686 44732 686 44760
rect -686 43708 602 44732
rect 666 43708 686 44732
rect -686 43680 686 43708
rect -686 43412 686 43440
rect -686 42388 602 43412
rect 666 42388 686 43412
rect -686 42360 686 42388
rect -686 42092 686 42120
rect -686 41068 602 42092
rect 666 41068 686 42092
rect -686 41040 686 41068
rect -686 40772 686 40800
rect -686 39748 602 40772
rect 666 39748 686 40772
rect -686 39720 686 39748
rect -686 39452 686 39480
rect -686 38428 602 39452
rect 666 38428 686 39452
rect -686 38400 686 38428
rect -686 38132 686 38160
rect -686 37108 602 38132
rect 666 37108 686 38132
rect -686 37080 686 37108
rect -686 36812 686 36840
rect -686 35788 602 36812
rect 666 35788 686 36812
rect -686 35760 686 35788
rect -686 35492 686 35520
rect -686 34468 602 35492
rect 666 34468 686 35492
rect -686 34440 686 34468
rect -686 34172 686 34200
rect -686 33148 602 34172
rect 666 33148 686 34172
rect -686 33120 686 33148
rect -686 32852 686 32880
rect -686 31828 602 32852
rect 666 31828 686 32852
rect -686 31800 686 31828
rect -686 31532 686 31560
rect -686 30508 602 31532
rect 666 30508 686 31532
rect -686 30480 686 30508
rect -686 30212 686 30240
rect -686 29188 602 30212
rect 666 29188 686 30212
rect -686 29160 686 29188
rect -686 28892 686 28920
rect -686 27868 602 28892
rect 666 27868 686 28892
rect -686 27840 686 27868
rect -686 27572 686 27600
rect -686 26548 602 27572
rect 666 26548 686 27572
rect -686 26520 686 26548
rect -686 26252 686 26280
rect -686 25228 602 26252
rect 666 25228 686 26252
rect -686 25200 686 25228
rect -686 24932 686 24960
rect -686 23908 602 24932
rect 666 23908 686 24932
rect -686 23880 686 23908
rect -686 23612 686 23640
rect -686 22588 602 23612
rect 666 22588 686 23612
rect -686 22560 686 22588
rect -686 22292 686 22320
rect -686 21268 602 22292
rect 666 21268 686 22292
rect -686 21240 686 21268
rect -686 20972 686 21000
rect -686 19948 602 20972
rect 666 19948 686 20972
rect -686 19920 686 19948
rect -686 19652 686 19680
rect -686 18628 602 19652
rect 666 18628 686 19652
rect -686 18600 686 18628
rect -686 18332 686 18360
rect -686 17308 602 18332
rect 666 17308 686 18332
rect -686 17280 686 17308
rect -686 17012 686 17040
rect -686 15988 602 17012
rect 666 15988 686 17012
rect -686 15960 686 15988
rect -686 15692 686 15720
rect -686 14668 602 15692
rect 666 14668 686 15692
rect -686 14640 686 14668
rect -686 14372 686 14400
rect -686 13348 602 14372
rect 666 13348 686 14372
rect -686 13320 686 13348
rect -686 13052 686 13080
rect -686 12028 602 13052
rect 666 12028 686 13052
rect -686 12000 686 12028
rect -686 11732 686 11760
rect -686 10708 602 11732
rect 666 10708 686 11732
rect -686 10680 686 10708
rect -686 10412 686 10440
rect -686 9388 602 10412
rect 666 9388 686 10412
rect -686 9360 686 9388
rect -686 9092 686 9120
rect -686 8068 602 9092
rect 666 8068 686 9092
rect -686 8040 686 8068
rect -686 7772 686 7800
rect -686 6748 602 7772
rect 666 6748 686 7772
rect -686 6720 686 6748
rect -686 6452 686 6480
rect -686 5428 602 6452
rect 666 5428 686 6452
rect -686 5400 686 5428
rect -686 5132 686 5160
rect -686 4108 602 5132
rect 666 4108 686 5132
rect -686 4080 686 4108
rect -686 3812 686 3840
rect -686 2788 602 3812
rect 666 2788 686 3812
rect -686 2760 686 2788
rect -686 2492 686 2520
rect -686 1468 602 2492
rect 666 1468 686 2492
rect -686 1440 686 1468
rect -686 1172 686 1200
rect -686 148 602 1172
rect 666 148 686 1172
rect -686 120 686 148
rect -686 -148 686 -120
rect -686 -1172 602 -148
rect 666 -1172 686 -148
rect -686 -1200 686 -1172
rect -686 -1468 686 -1440
rect -686 -2492 602 -1468
rect 666 -2492 686 -1468
rect -686 -2520 686 -2492
rect -686 -2788 686 -2760
rect -686 -3812 602 -2788
rect 666 -3812 686 -2788
rect -686 -3840 686 -3812
rect -686 -4108 686 -4080
rect -686 -5132 602 -4108
rect 666 -5132 686 -4108
rect -686 -5160 686 -5132
rect -686 -5428 686 -5400
rect -686 -6452 602 -5428
rect 666 -6452 686 -5428
rect -686 -6480 686 -6452
rect -686 -6748 686 -6720
rect -686 -7772 602 -6748
rect 666 -7772 686 -6748
rect -686 -7800 686 -7772
rect -686 -8068 686 -8040
rect -686 -9092 602 -8068
rect 666 -9092 686 -8068
rect -686 -9120 686 -9092
rect -686 -9388 686 -9360
rect -686 -10412 602 -9388
rect 666 -10412 686 -9388
rect -686 -10440 686 -10412
rect -686 -10708 686 -10680
rect -686 -11732 602 -10708
rect 666 -11732 686 -10708
rect -686 -11760 686 -11732
rect -686 -12028 686 -12000
rect -686 -13052 602 -12028
rect 666 -13052 686 -12028
rect -686 -13080 686 -13052
rect -686 -13348 686 -13320
rect -686 -14372 602 -13348
rect 666 -14372 686 -13348
rect -686 -14400 686 -14372
rect -686 -14668 686 -14640
rect -686 -15692 602 -14668
rect 666 -15692 686 -14668
rect -686 -15720 686 -15692
rect -686 -15988 686 -15960
rect -686 -17012 602 -15988
rect 666 -17012 686 -15988
rect -686 -17040 686 -17012
rect -686 -17308 686 -17280
rect -686 -18332 602 -17308
rect 666 -18332 686 -17308
rect -686 -18360 686 -18332
rect -686 -18628 686 -18600
rect -686 -19652 602 -18628
rect 666 -19652 686 -18628
rect -686 -19680 686 -19652
rect -686 -19948 686 -19920
rect -686 -20972 602 -19948
rect 666 -20972 686 -19948
rect -686 -21000 686 -20972
rect -686 -21268 686 -21240
rect -686 -22292 602 -21268
rect 666 -22292 686 -21268
rect -686 -22320 686 -22292
rect -686 -22588 686 -22560
rect -686 -23612 602 -22588
rect 666 -23612 686 -22588
rect -686 -23640 686 -23612
rect -686 -23908 686 -23880
rect -686 -24932 602 -23908
rect 666 -24932 686 -23908
rect -686 -24960 686 -24932
rect -686 -25228 686 -25200
rect -686 -26252 602 -25228
rect 666 -26252 686 -25228
rect -686 -26280 686 -26252
rect -686 -26548 686 -26520
rect -686 -27572 602 -26548
rect 666 -27572 686 -26548
rect -686 -27600 686 -27572
rect -686 -27868 686 -27840
rect -686 -28892 602 -27868
rect 666 -28892 686 -27868
rect -686 -28920 686 -28892
rect -686 -29188 686 -29160
rect -686 -30212 602 -29188
rect 666 -30212 686 -29188
rect -686 -30240 686 -30212
rect -686 -30508 686 -30480
rect -686 -31532 602 -30508
rect 666 -31532 686 -30508
rect -686 -31560 686 -31532
rect -686 -31828 686 -31800
rect -686 -32852 602 -31828
rect 666 -32852 686 -31828
rect -686 -32880 686 -32852
rect -686 -33148 686 -33120
rect -686 -34172 602 -33148
rect 666 -34172 686 -33148
rect -686 -34200 686 -34172
rect -686 -34468 686 -34440
rect -686 -35492 602 -34468
rect 666 -35492 686 -34468
rect -686 -35520 686 -35492
rect -686 -35788 686 -35760
rect -686 -36812 602 -35788
rect 666 -36812 686 -35788
rect -686 -36840 686 -36812
rect -686 -37108 686 -37080
rect -686 -38132 602 -37108
rect 666 -38132 686 -37108
rect -686 -38160 686 -38132
rect -686 -38428 686 -38400
rect -686 -39452 602 -38428
rect 666 -39452 686 -38428
rect -686 -39480 686 -39452
rect -686 -39748 686 -39720
rect -686 -40772 602 -39748
rect 666 -40772 686 -39748
rect -686 -40800 686 -40772
rect -686 -41068 686 -41040
rect -686 -42092 602 -41068
rect 666 -42092 686 -41068
rect -686 -42120 686 -42092
rect -686 -42388 686 -42360
rect -686 -43412 602 -42388
rect 666 -43412 686 -42388
rect -686 -43440 686 -43412
rect -686 -43708 686 -43680
rect -686 -44732 602 -43708
rect 666 -44732 686 -43708
rect -686 -44760 686 -44732
rect -686 -45028 686 -45000
rect -686 -46052 602 -45028
rect 666 -46052 686 -45028
rect -686 -46080 686 -46052
rect -686 -46348 686 -46320
rect -686 -47372 602 -46348
rect 666 -47372 686 -46348
rect -686 -47400 686 -47372
rect -686 -47668 686 -47640
rect -686 -48692 602 -47668
rect 666 -48692 686 -47668
rect -686 -48720 686 -48692
rect -686 -48988 686 -48960
rect -686 -50012 602 -48988
rect 666 -50012 686 -48988
rect -686 -50040 686 -50012
rect -686 -50308 686 -50280
rect -686 -51332 602 -50308
rect 666 -51332 686 -50308
rect -686 -51360 686 -51332
rect -686 -51628 686 -51600
rect -686 -52652 602 -51628
rect 666 -52652 686 -51628
rect -686 -52680 686 -52652
rect -686 -52948 686 -52920
rect -686 -53972 602 -52948
rect 666 -53972 686 -52948
rect -686 -54000 686 -53972
rect -686 -54268 686 -54240
rect -686 -55292 602 -54268
rect 666 -55292 686 -54268
rect -686 -55320 686 -55292
rect -686 -55588 686 -55560
rect -686 -56612 602 -55588
rect 666 -56612 686 -55588
rect -686 -56640 686 -56612
rect -686 -56908 686 -56880
rect -686 -57932 602 -56908
rect 666 -57932 686 -56908
rect -686 -57960 686 -57932
rect -686 -58228 686 -58200
rect -686 -59252 602 -58228
rect 666 -59252 686 -58228
rect -686 -59280 686 -59252
rect -686 -59548 686 -59520
rect -686 -60572 602 -59548
rect 666 -60572 686 -59548
rect -686 -60600 686 -60572
rect -686 -60868 686 -60840
rect -686 -61892 602 -60868
rect 666 -61892 686 -60868
rect -686 -61920 686 -61892
rect -686 -62188 686 -62160
rect -686 -63212 602 -62188
rect 666 -63212 686 -62188
rect -686 -63240 686 -63212
rect -686 -63508 686 -63480
rect -686 -64532 602 -63508
rect 666 -64532 686 -63508
rect -686 -64560 686 -64532
rect -686 -64828 686 -64800
rect -686 -65852 602 -64828
rect 666 -65852 686 -64828
rect -686 -65880 686 -65852
rect -686 -66148 686 -66120
rect -686 -67172 602 -66148
rect 666 -67172 686 -66148
rect -686 -67200 686 -67172
rect -686 -67468 686 -67440
rect -686 -68492 602 -67468
rect 666 -68492 686 -67468
rect -686 -68520 686 -68492
rect -686 -68788 686 -68760
rect -686 -69812 602 -68788
rect 666 -69812 686 -68788
rect -686 -69840 686 -69812
rect -686 -70108 686 -70080
rect -686 -71132 602 -70108
rect 666 -71132 686 -70108
rect -686 -71160 686 -71132
rect -686 -71428 686 -71400
rect -686 -72452 602 -71428
rect 666 -72452 686 -71428
rect -686 -72480 686 -72452
rect -686 -72748 686 -72720
rect -686 -73772 602 -72748
rect 666 -73772 686 -72748
rect -686 -73800 686 -73772
rect -686 -74068 686 -74040
rect -686 -75092 602 -74068
rect 666 -75092 686 -74068
rect -686 -75120 686 -75092
rect -686 -75388 686 -75360
rect -686 -76412 602 -75388
rect 666 -76412 686 -75388
rect -686 -76440 686 -76412
rect -686 -76708 686 -76680
rect -686 -77732 602 -76708
rect 666 -77732 686 -76708
rect -686 -77760 686 -77732
rect -686 -78028 686 -78000
rect -686 -79052 602 -78028
rect 666 -79052 686 -78028
rect -686 -79080 686 -79052
rect -686 -79348 686 -79320
rect -686 -80372 602 -79348
rect 666 -80372 686 -79348
rect -686 -80400 686 -80372
rect -686 -80668 686 -80640
rect -686 -81692 602 -80668
rect 666 -81692 686 -80668
rect -686 -81720 686 -81692
rect -686 -81988 686 -81960
rect -686 -83012 602 -81988
rect 666 -83012 686 -81988
rect -686 -83040 686 -83012
rect -686 -83308 686 -83280
rect -686 -84332 602 -83308
rect 666 -84332 686 -83308
rect -686 -84360 686 -84332
<< via3 >>
rect 602 83308 666 84332
rect 602 81988 666 83012
rect 602 80668 666 81692
rect 602 79348 666 80372
rect 602 78028 666 79052
rect 602 76708 666 77732
rect 602 75388 666 76412
rect 602 74068 666 75092
rect 602 72748 666 73772
rect 602 71428 666 72452
rect 602 70108 666 71132
rect 602 68788 666 69812
rect 602 67468 666 68492
rect 602 66148 666 67172
rect 602 64828 666 65852
rect 602 63508 666 64532
rect 602 62188 666 63212
rect 602 60868 666 61892
rect 602 59548 666 60572
rect 602 58228 666 59252
rect 602 56908 666 57932
rect 602 55588 666 56612
rect 602 54268 666 55292
rect 602 52948 666 53972
rect 602 51628 666 52652
rect 602 50308 666 51332
rect 602 48988 666 50012
rect 602 47668 666 48692
rect 602 46348 666 47372
rect 602 45028 666 46052
rect 602 43708 666 44732
rect 602 42388 666 43412
rect 602 41068 666 42092
rect 602 39748 666 40772
rect 602 38428 666 39452
rect 602 37108 666 38132
rect 602 35788 666 36812
rect 602 34468 666 35492
rect 602 33148 666 34172
rect 602 31828 666 32852
rect 602 30508 666 31532
rect 602 29188 666 30212
rect 602 27868 666 28892
rect 602 26548 666 27572
rect 602 25228 666 26252
rect 602 23908 666 24932
rect 602 22588 666 23612
rect 602 21268 666 22292
rect 602 19948 666 20972
rect 602 18628 666 19652
rect 602 17308 666 18332
rect 602 15988 666 17012
rect 602 14668 666 15692
rect 602 13348 666 14372
rect 602 12028 666 13052
rect 602 10708 666 11732
rect 602 9388 666 10412
rect 602 8068 666 9092
rect 602 6748 666 7772
rect 602 5428 666 6452
rect 602 4108 666 5132
rect 602 2788 666 3812
rect 602 1468 666 2492
rect 602 148 666 1172
rect 602 -1172 666 -148
rect 602 -2492 666 -1468
rect 602 -3812 666 -2788
rect 602 -5132 666 -4108
rect 602 -6452 666 -5428
rect 602 -7772 666 -6748
rect 602 -9092 666 -8068
rect 602 -10412 666 -9388
rect 602 -11732 666 -10708
rect 602 -13052 666 -12028
rect 602 -14372 666 -13348
rect 602 -15692 666 -14668
rect 602 -17012 666 -15988
rect 602 -18332 666 -17308
rect 602 -19652 666 -18628
rect 602 -20972 666 -19948
rect 602 -22292 666 -21268
rect 602 -23612 666 -22588
rect 602 -24932 666 -23908
rect 602 -26252 666 -25228
rect 602 -27572 666 -26548
rect 602 -28892 666 -27868
rect 602 -30212 666 -29188
rect 602 -31532 666 -30508
rect 602 -32852 666 -31828
rect 602 -34172 666 -33148
rect 602 -35492 666 -34468
rect 602 -36812 666 -35788
rect 602 -38132 666 -37108
rect 602 -39452 666 -38428
rect 602 -40772 666 -39748
rect 602 -42092 666 -41068
rect 602 -43412 666 -42388
rect 602 -44732 666 -43708
rect 602 -46052 666 -45028
rect 602 -47372 666 -46348
rect 602 -48692 666 -47668
rect 602 -50012 666 -48988
rect 602 -51332 666 -50308
rect 602 -52652 666 -51628
rect 602 -53972 666 -52948
rect 602 -55292 666 -54268
rect 602 -56612 666 -55588
rect 602 -57932 666 -56908
rect 602 -59252 666 -58228
rect 602 -60572 666 -59548
rect 602 -61892 666 -60868
rect 602 -63212 666 -62188
rect 602 -64532 666 -63508
rect 602 -65852 666 -64828
rect 602 -67172 666 -66148
rect 602 -68492 666 -67468
rect 602 -69812 666 -68788
rect 602 -71132 666 -70108
rect 602 -72452 666 -71428
rect 602 -73772 666 -72748
rect 602 -75092 666 -74068
rect 602 -76412 666 -75388
rect 602 -77732 666 -76708
rect 602 -79052 666 -78028
rect 602 -80372 666 -79348
rect 602 -81692 666 -80668
rect 602 -83012 666 -81988
rect 602 -84332 666 -83308
<< mimcap >>
rect -646 84280 354 84320
rect -646 83360 -606 84280
rect 314 83360 354 84280
rect -646 83320 354 83360
rect -646 82960 354 83000
rect -646 82040 -606 82960
rect 314 82040 354 82960
rect -646 82000 354 82040
rect -646 81640 354 81680
rect -646 80720 -606 81640
rect 314 80720 354 81640
rect -646 80680 354 80720
rect -646 80320 354 80360
rect -646 79400 -606 80320
rect 314 79400 354 80320
rect -646 79360 354 79400
rect -646 79000 354 79040
rect -646 78080 -606 79000
rect 314 78080 354 79000
rect -646 78040 354 78080
rect -646 77680 354 77720
rect -646 76760 -606 77680
rect 314 76760 354 77680
rect -646 76720 354 76760
rect -646 76360 354 76400
rect -646 75440 -606 76360
rect 314 75440 354 76360
rect -646 75400 354 75440
rect -646 75040 354 75080
rect -646 74120 -606 75040
rect 314 74120 354 75040
rect -646 74080 354 74120
rect -646 73720 354 73760
rect -646 72800 -606 73720
rect 314 72800 354 73720
rect -646 72760 354 72800
rect -646 72400 354 72440
rect -646 71480 -606 72400
rect 314 71480 354 72400
rect -646 71440 354 71480
rect -646 71080 354 71120
rect -646 70160 -606 71080
rect 314 70160 354 71080
rect -646 70120 354 70160
rect -646 69760 354 69800
rect -646 68840 -606 69760
rect 314 68840 354 69760
rect -646 68800 354 68840
rect -646 68440 354 68480
rect -646 67520 -606 68440
rect 314 67520 354 68440
rect -646 67480 354 67520
rect -646 67120 354 67160
rect -646 66200 -606 67120
rect 314 66200 354 67120
rect -646 66160 354 66200
rect -646 65800 354 65840
rect -646 64880 -606 65800
rect 314 64880 354 65800
rect -646 64840 354 64880
rect -646 64480 354 64520
rect -646 63560 -606 64480
rect 314 63560 354 64480
rect -646 63520 354 63560
rect -646 63160 354 63200
rect -646 62240 -606 63160
rect 314 62240 354 63160
rect -646 62200 354 62240
rect -646 61840 354 61880
rect -646 60920 -606 61840
rect 314 60920 354 61840
rect -646 60880 354 60920
rect -646 60520 354 60560
rect -646 59600 -606 60520
rect 314 59600 354 60520
rect -646 59560 354 59600
rect -646 59200 354 59240
rect -646 58280 -606 59200
rect 314 58280 354 59200
rect -646 58240 354 58280
rect -646 57880 354 57920
rect -646 56960 -606 57880
rect 314 56960 354 57880
rect -646 56920 354 56960
rect -646 56560 354 56600
rect -646 55640 -606 56560
rect 314 55640 354 56560
rect -646 55600 354 55640
rect -646 55240 354 55280
rect -646 54320 -606 55240
rect 314 54320 354 55240
rect -646 54280 354 54320
rect -646 53920 354 53960
rect -646 53000 -606 53920
rect 314 53000 354 53920
rect -646 52960 354 53000
rect -646 52600 354 52640
rect -646 51680 -606 52600
rect 314 51680 354 52600
rect -646 51640 354 51680
rect -646 51280 354 51320
rect -646 50360 -606 51280
rect 314 50360 354 51280
rect -646 50320 354 50360
rect -646 49960 354 50000
rect -646 49040 -606 49960
rect 314 49040 354 49960
rect -646 49000 354 49040
rect -646 48640 354 48680
rect -646 47720 -606 48640
rect 314 47720 354 48640
rect -646 47680 354 47720
rect -646 47320 354 47360
rect -646 46400 -606 47320
rect 314 46400 354 47320
rect -646 46360 354 46400
rect -646 46000 354 46040
rect -646 45080 -606 46000
rect 314 45080 354 46000
rect -646 45040 354 45080
rect -646 44680 354 44720
rect -646 43760 -606 44680
rect 314 43760 354 44680
rect -646 43720 354 43760
rect -646 43360 354 43400
rect -646 42440 -606 43360
rect 314 42440 354 43360
rect -646 42400 354 42440
rect -646 42040 354 42080
rect -646 41120 -606 42040
rect 314 41120 354 42040
rect -646 41080 354 41120
rect -646 40720 354 40760
rect -646 39800 -606 40720
rect 314 39800 354 40720
rect -646 39760 354 39800
rect -646 39400 354 39440
rect -646 38480 -606 39400
rect 314 38480 354 39400
rect -646 38440 354 38480
rect -646 38080 354 38120
rect -646 37160 -606 38080
rect 314 37160 354 38080
rect -646 37120 354 37160
rect -646 36760 354 36800
rect -646 35840 -606 36760
rect 314 35840 354 36760
rect -646 35800 354 35840
rect -646 35440 354 35480
rect -646 34520 -606 35440
rect 314 34520 354 35440
rect -646 34480 354 34520
rect -646 34120 354 34160
rect -646 33200 -606 34120
rect 314 33200 354 34120
rect -646 33160 354 33200
rect -646 32800 354 32840
rect -646 31880 -606 32800
rect 314 31880 354 32800
rect -646 31840 354 31880
rect -646 31480 354 31520
rect -646 30560 -606 31480
rect 314 30560 354 31480
rect -646 30520 354 30560
rect -646 30160 354 30200
rect -646 29240 -606 30160
rect 314 29240 354 30160
rect -646 29200 354 29240
rect -646 28840 354 28880
rect -646 27920 -606 28840
rect 314 27920 354 28840
rect -646 27880 354 27920
rect -646 27520 354 27560
rect -646 26600 -606 27520
rect 314 26600 354 27520
rect -646 26560 354 26600
rect -646 26200 354 26240
rect -646 25280 -606 26200
rect 314 25280 354 26200
rect -646 25240 354 25280
rect -646 24880 354 24920
rect -646 23960 -606 24880
rect 314 23960 354 24880
rect -646 23920 354 23960
rect -646 23560 354 23600
rect -646 22640 -606 23560
rect 314 22640 354 23560
rect -646 22600 354 22640
rect -646 22240 354 22280
rect -646 21320 -606 22240
rect 314 21320 354 22240
rect -646 21280 354 21320
rect -646 20920 354 20960
rect -646 20000 -606 20920
rect 314 20000 354 20920
rect -646 19960 354 20000
rect -646 19600 354 19640
rect -646 18680 -606 19600
rect 314 18680 354 19600
rect -646 18640 354 18680
rect -646 18280 354 18320
rect -646 17360 -606 18280
rect 314 17360 354 18280
rect -646 17320 354 17360
rect -646 16960 354 17000
rect -646 16040 -606 16960
rect 314 16040 354 16960
rect -646 16000 354 16040
rect -646 15640 354 15680
rect -646 14720 -606 15640
rect 314 14720 354 15640
rect -646 14680 354 14720
rect -646 14320 354 14360
rect -646 13400 -606 14320
rect 314 13400 354 14320
rect -646 13360 354 13400
rect -646 13000 354 13040
rect -646 12080 -606 13000
rect 314 12080 354 13000
rect -646 12040 354 12080
rect -646 11680 354 11720
rect -646 10760 -606 11680
rect 314 10760 354 11680
rect -646 10720 354 10760
rect -646 10360 354 10400
rect -646 9440 -606 10360
rect 314 9440 354 10360
rect -646 9400 354 9440
rect -646 9040 354 9080
rect -646 8120 -606 9040
rect 314 8120 354 9040
rect -646 8080 354 8120
rect -646 7720 354 7760
rect -646 6800 -606 7720
rect 314 6800 354 7720
rect -646 6760 354 6800
rect -646 6400 354 6440
rect -646 5480 -606 6400
rect 314 5480 354 6400
rect -646 5440 354 5480
rect -646 5080 354 5120
rect -646 4160 -606 5080
rect 314 4160 354 5080
rect -646 4120 354 4160
rect -646 3760 354 3800
rect -646 2840 -606 3760
rect 314 2840 354 3760
rect -646 2800 354 2840
rect -646 2440 354 2480
rect -646 1520 -606 2440
rect 314 1520 354 2440
rect -646 1480 354 1520
rect -646 1120 354 1160
rect -646 200 -606 1120
rect 314 200 354 1120
rect -646 160 354 200
rect -646 -200 354 -160
rect -646 -1120 -606 -200
rect 314 -1120 354 -200
rect -646 -1160 354 -1120
rect -646 -1520 354 -1480
rect -646 -2440 -606 -1520
rect 314 -2440 354 -1520
rect -646 -2480 354 -2440
rect -646 -2840 354 -2800
rect -646 -3760 -606 -2840
rect 314 -3760 354 -2840
rect -646 -3800 354 -3760
rect -646 -4160 354 -4120
rect -646 -5080 -606 -4160
rect 314 -5080 354 -4160
rect -646 -5120 354 -5080
rect -646 -5480 354 -5440
rect -646 -6400 -606 -5480
rect 314 -6400 354 -5480
rect -646 -6440 354 -6400
rect -646 -6800 354 -6760
rect -646 -7720 -606 -6800
rect 314 -7720 354 -6800
rect -646 -7760 354 -7720
rect -646 -8120 354 -8080
rect -646 -9040 -606 -8120
rect 314 -9040 354 -8120
rect -646 -9080 354 -9040
rect -646 -9440 354 -9400
rect -646 -10360 -606 -9440
rect 314 -10360 354 -9440
rect -646 -10400 354 -10360
rect -646 -10760 354 -10720
rect -646 -11680 -606 -10760
rect 314 -11680 354 -10760
rect -646 -11720 354 -11680
rect -646 -12080 354 -12040
rect -646 -13000 -606 -12080
rect 314 -13000 354 -12080
rect -646 -13040 354 -13000
rect -646 -13400 354 -13360
rect -646 -14320 -606 -13400
rect 314 -14320 354 -13400
rect -646 -14360 354 -14320
rect -646 -14720 354 -14680
rect -646 -15640 -606 -14720
rect 314 -15640 354 -14720
rect -646 -15680 354 -15640
rect -646 -16040 354 -16000
rect -646 -16960 -606 -16040
rect 314 -16960 354 -16040
rect -646 -17000 354 -16960
rect -646 -17360 354 -17320
rect -646 -18280 -606 -17360
rect 314 -18280 354 -17360
rect -646 -18320 354 -18280
rect -646 -18680 354 -18640
rect -646 -19600 -606 -18680
rect 314 -19600 354 -18680
rect -646 -19640 354 -19600
rect -646 -20000 354 -19960
rect -646 -20920 -606 -20000
rect 314 -20920 354 -20000
rect -646 -20960 354 -20920
rect -646 -21320 354 -21280
rect -646 -22240 -606 -21320
rect 314 -22240 354 -21320
rect -646 -22280 354 -22240
rect -646 -22640 354 -22600
rect -646 -23560 -606 -22640
rect 314 -23560 354 -22640
rect -646 -23600 354 -23560
rect -646 -23960 354 -23920
rect -646 -24880 -606 -23960
rect 314 -24880 354 -23960
rect -646 -24920 354 -24880
rect -646 -25280 354 -25240
rect -646 -26200 -606 -25280
rect 314 -26200 354 -25280
rect -646 -26240 354 -26200
rect -646 -26600 354 -26560
rect -646 -27520 -606 -26600
rect 314 -27520 354 -26600
rect -646 -27560 354 -27520
rect -646 -27920 354 -27880
rect -646 -28840 -606 -27920
rect 314 -28840 354 -27920
rect -646 -28880 354 -28840
rect -646 -29240 354 -29200
rect -646 -30160 -606 -29240
rect 314 -30160 354 -29240
rect -646 -30200 354 -30160
rect -646 -30560 354 -30520
rect -646 -31480 -606 -30560
rect 314 -31480 354 -30560
rect -646 -31520 354 -31480
rect -646 -31880 354 -31840
rect -646 -32800 -606 -31880
rect 314 -32800 354 -31880
rect -646 -32840 354 -32800
rect -646 -33200 354 -33160
rect -646 -34120 -606 -33200
rect 314 -34120 354 -33200
rect -646 -34160 354 -34120
rect -646 -34520 354 -34480
rect -646 -35440 -606 -34520
rect 314 -35440 354 -34520
rect -646 -35480 354 -35440
rect -646 -35840 354 -35800
rect -646 -36760 -606 -35840
rect 314 -36760 354 -35840
rect -646 -36800 354 -36760
rect -646 -37160 354 -37120
rect -646 -38080 -606 -37160
rect 314 -38080 354 -37160
rect -646 -38120 354 -38080
rect -646 -38480 354 -38440
rect -646 -39400 -606 -38480
rect 314 -39400 354 -38480
rect -646 -39440 354 -39400
rect -646 -39800 354 -39760
rect -646 -40720 -606 -39800
rect 314 -40720 354 -39800
rect -646 -40760 354 -40720
rect -646 -41120 354 -41080
rect -646 -42040 -606 -41120
rect 314 -42040 354 -41120
rect -646 -42080 354 -42040
rect -646 -42440 354 -42400
rect -646 -43360 -606 -42440
rect 314 -43360 354 -42440
rect -646 -43400 354 -43360
rect -646 -43760 354 -43720
rect -646 -44680 -606 -43760
rect 314 -44680 354 -43760
rect -646 -44720 354 -44680
rect -646 -45080 354 -45040
rect -646 -46000 -606 -45080
rect 314 -46000 354 -45080
rect -646 -46040 354 -46000
rect -646 -46400 354 -46360
rect -646 -47320 -606 -46400
rect 314 -47320 354 -46400
rect -646 -47360 354 -47320
rect -646 -47720 354 -47680
rect -646 -48640 -606 -47720
rect 314 -48640 354 -47720
rect -646 -48680 354 -48640
rect -646 -49040 354 -49000
rect -646 -49960 -606 -49040
rect 314 -49960 354 -49040
rect -646 -50000 354 -49960
rect -646 -50360 354 -50320
rect -646 -51280 -606 -50360
rect 314 -51280 354 -50360
rect -646 -51320 354 -51280
rect -646 -51680 354 -51640
rect -646 -52600 -606 -51680
rect 314 -52600 354 -51680
rect -646 -52640 354 -52600
rect -646 -53000 354 -52960
rect -646 -53920 -606 -53000
rect 314 -53920 354 -53000
rect -646 -53960 354 -53920
rect -646 -54320 354 -54280
rect -646 -55240 -606 -54320
rect 314 -55240 354 -54320
rect -646 -55280 354 -55240
rect -646 -55640 354 -55600
rect -646 -56560 -606 -55640
rect 314 -56560 354 -55640
rect -646 -56600 354 -56560
rect -646 -56960 354 -56920
rect -646 -57880 -606 -56960
rect 314 -57880 354 -56960
rect -646 -57920 354 -57880
rect -646 -58280 354 -58240
rect -646 -59200 -606 -58280
rect 314 -59200 354 -58280
rect -646 -59240 354 -59200
rect -646 -59600 354 -59560
rect -646 -60520 -606 -59600
rect 314 -60520 354 -59600
rect -646 -60560 354 -60520
rect -646 -60920 354 -60880
rect -646 -61840 -606 -60920
rect 314 -61840 354 -60920
rect -646 -61880 354 -61840
rect -646 -62240 354 -62200
rect -646 -63160 -606 -62240
rect 314 -63160 354 -62240
rect -646 -63200 354 -63160
rect -646 -63560 354 -63520
rect -646 -64480 -606 -63560
rect 314 -64480 354 -63560
rect -646 -64520 354 -64480
rect -646 -64880 354 -64840
rect -646 -65800 -606 -64880
rect 314 -65800 354 -64880
rect -646 -65840 354 -65800
rect -646 -66200 354 -66160
rect -646 -67120 -606 -66200
rect 314 -67120 354 -66200
rect -646 -67160 354 -67120
rect -646 -67520 354 -67480
rect -646 -68440 -606 -67520
rect 314 -68440 354 -67520
rect -646 -68480 354 -68440
rect -646 -68840 354 -68800
rect -646 -69760 -606 -68840
rect 314 -69760 354 -68840
rect -646 -69800 354 -69760
rect -646 -70160 354 -70120
rect -646 -71080 -606 -70160
rect 314 -71080 354 -70160
rect -646 -71120 354 -71080
rect -646 -71480 354 -71440
rect -646 -72400 -606 -71480
rect 314 -72400 354 -71480
rect -646 -72440 354 -72400
rect -646 -72800 354 -72760
rect -646 -73720 -606 -72800
rect 314 -73720 354 -72800
rect -646 -73760 354 -73720
rect -646 -74120 354 -74080
rect -646 -75040 -606 -74120
rect 314 -75040 354 -74120
rect -646 -75080 354 -75040
rect -646 -75440 354 -75400
rect -646 -76360 -606 -75440
rect 314 -76360 354 -75440
rect -646 -76400 354 -76360
rect -646 -76760 354 -76720
rect -646 -77680 -606 -76760
rect 314 -77680 354 -76760
rect -646 -77720 354 -77680
rect -646 -78080 354 -78040
rect -646 -79000 -606 -78080
rect 314 -79000 354 -78080
rect -646 -79040 354 -79000
rect -646 -79400 354 -79360
rect -646 -80320 -606 -79400
rect 314 -80320 354 -79400
rect -646 -80360 354 -80320
rect -646 -80720 354 -80680
rect -646 -81640 -606 -80720
rect 314 -81640 354 -80720
rect -646 -81680 354 -81640
rect -646 -82040 354 -82000
rect -646 -82960 -606 -82040
rect 314 -82960 354 -82040
rect -646 -83000 354 -82960
rect -646 -83360 354 -83320
rect -646 -84280 -606 -83360
rect 314 -84280 354 -83360
rect -646 -84320 354 -84280
<< mimcapcontact >>
rect -606 83360 314 84280
rect -606 82040 314 82960
rect -606 80720 314 81640
rect -606 79400 314 80320
rect -606 78080 314 79000
rect -606 76760 314 77680
rect -606 75440 314 76360
rect -606 74120 314 75040
rect -606 72800 314 73720
rect -606 71480 314 72400
rect -606 70160 314 71080
rect -606 68840 314 69760
rect -606 67520 314 68440
rect -606 66200 314 67120
rect -606 64880 314 65800
rect -606 63560 314 64480
rect -606 62240 314 63160
rect -606 60920 314 61840
rect -606 59600 314 60520
rect -606 58280 314 59200
rect -606 56960 314 57880
rect -606 55640 314 56560
rect -606 54320 314 55240
rect -606 53000 314 53920
rect -606 51680 314 52600
rect -606 50360 314 51280
rect -606 49040 314 49960
rect -606 47720 314 48640
rect -606 46400 314 47320
rect -606 45080 314 46000
rect -606 43760 314 44680
rect -606 42440 314 43360
rect -606 41120 314 42040
rect -606 39800 314 40720
rect -606 38480 314 39400
rect -606 37160 314 38080
rect -606 35840 314 36760
rect -606 34520 314 35440
rect -606 33200 314 34120
rect -606 31880 314 32800
rect -606 30560 314 31480
rect -606 29240 314 30160
rect -606 27920 314 28840
rect -606 26600 314 27520
rect -606 25280 314 26200
rect -606 23960 314 24880
rect -606 22640 314 23560
rect -606 21320 314 22240
rect -606 20000 314 20920
rect -606 18680 314 19600
rect -606 17360 314 18280
rect -606 16040 314 16960
rect -606 14720 314 15640
rect -606 13400 314 14320
rect -606 12080 314 13000
rect -606 10760 314 11680
rect -606 9440 314 10360
rect -606 8120 314 9040
rect -606 6800 314 7720
rect -606 5480 314 6400
rect -606 4160 314 5080
rect -606 2840 314 3760
rect -606 1520 314 2440
rect -606 200 314 1120
rect -606 -1120 314 -200
rect -606 -2440 314 -1520
rect -606 -3760 314 -2840
rect -606 -5080 314 -4160
rect -606 -6400 314 -5480
rect -606 -7720 314 -6800
rect -606 -9040 314 -8120
rect -606 -10360 314 -9440
rect -606 -11680 314 -10760
rect -606 -13000 314 -12080
rect -606 -14320 314 -13400
rect -606 -15640 314 -14720
rect -606 -16960 314 -16040
rect -606 -18280 314 -17360
rect -606 -19600 314 -18680
rect -606 -20920 314 -20000
rect -606 -22240 314 -21320
rect -606 -23560 314 -22640
rect -606 -24880 314 -23960
rect -606 -26200 314 -25280
rect -606 -27520 314 -26600
rect -606 -28840 314 -27920
rect -606 -30160 314 -29240
rect -606 -31480 314 -30560
rect -606 -32800 314 -31880
rect -606 -34120 314 -33200
rect -606 -35440 314 -34520
rect -606 -36760 314 -35840
rect -606 -38080 314 -37160
rect -606 -39400 314 -38480
rect -606 -40720 314 -39800
rect -606 -42040 314 -41120
rect -606 -43360 314 -42440
rect -606 -44680 314 -43760
rect -606 -46000 314 -45080
rect -606 -47320 314 -46400
rect -606 -48640 314 -47720
rect -606 -49960 314 -49040
rect -606 -51280 314 -50360
rect -606 -52600 314 -51680
rect -606 -53920 314 -53000
rect -606 -55240 314 -54320
rect -606 -56560 314 -55640
rect -606 -57880 314 -56960
rect -606 -59200 314 -58280
rect -606 -60520 314 -59600
rect -606 -61840 314 -60920
rect -606 -63160 314 -62240
rect -606 -64480 314 -63560
rect -606 -65800 314 -64880
rect -606 -67120 314 -66200
rect -606 -68440 314 -67520
rect -606 -69760 314 -68840
rect -606 -71080 314 -70160
rect -606 -72400 314 -71480
rect -606 -73720 314 -72800
rect -606 -75040 314 -74120
rect -606 -76360 314 -75440
rect -606 -77680 314 -76760
rect -606 -79000 314 -78080
rect -606 -80320 314 -79400
rect -606 -81640 314 -80720
rect -606 -82960 314 -82040
rect -606 -84280 314 -83360
<< metal4 >>
rect -198 84281 -94 84480
rect 582 84332 686 84480
rect -607 84280 315 84281
rect -607 83360 -606 84280
rect 314 83360 315 84280
rect -607 83359 315 83360
rect -198 82961 -94 83359
rect 582 83308 602 84332
rect 666 83308 686 84332
rect 582 83012 686 83308
rect -607 82960 315 82961
rect -607 82040 -606 82960
rect 314 82040 315 82960
rect -607 82039 315 82040
rect -198 81641 -94 82039
rect 582 81988 602 83012
rect 666 81988 686 83012
rect 582 81692 686 81988
rect -607 81640 315 81641
rect -607 80720 -606 81640
rect 314 80720 315 81640
rect -607 80719 315 80720
rect -198 80321 -94 80719
rect 582 80668 602 81692
rect 666 80668 686 81692
rect 582 80372 686 80668
rect -607 80320 315 80321
rect -607 79400 -606 80320
rect 314 79400 315 80320
rect -607 79399 315 79400
rect -198 79001 -94 79399
rect 582 79348 602 80372
rect 666 79348 686 80372
rect 582 79052 686 79348
rect -607 79000 315 79001
rect -607 78080 -606 79000
rect 314 78080 315 79000
rect -607 78079 315 78080
rect -198 77681 -94 78079
rect 582 78028 602 79052
rect 666 78028 686 79052
rect 582 77732 686 78028
rect -607 77680 315 77681
rect -607 76760 -606 77680
rect 314 76760 315 77680
rect -607 76759 315 76760
rect -198 76361 -94 76759
rect 582 76708 602 77732
rect 666 76708 686 77732
rect 582 76412 686 76708
rect -607 76360 315 76361
rect -607 75440 -606 76360
rect 314 75440 315 76360
rect -607 75439 315 75440
rect -198 75041 -94 75439
rect 582 75388 602 76412
rect 666 75388 686 76412
rect 582 75092 686 75388
rect -607 75040 315 75041
rect -607 74120 -606 75040
rect 314 74120 315 75040
rect -607 74119 315 74120
rect -198 73721 -94 74119
rect 582 74068 602 75092
rect 666 74068 686 75092
rect 582 73772 686 74068
rect -607 73720 315 73721
rect -607 72800 -606 73720
rect 314 72800 315 73720
rect -607 72799 315 72800
rect -198 72401 -94 72799
rect 582 72748 602 73772
rect 666 72748 686 73772
rect 582 72452 686 72748
rect -607 72400 315 72401
rect -607 71480 -606 72400
rect 314 71480 315 72400
rect -607 71479 315 71480
rect -198 71081 -94 71479
rect 582 71428 602 72452
rect 666 71428 686 72452
rect 582 71132 686 71428
rect -607 71080 315 71081
rect -607 70160 -606 71080
rect 314 70160 315 71080
rect -607 70159 315 70160
rect -198 69761 -94 70159
rect 582 70108 602 71132
rect 666 70108 686 71132
rect 582 69812 686 70108
rect -607 69760 315 69761
rect -607 68840 -606 69760
rect 314 68840 315 69760
rect -607 68839 315 68840
rect -198 68441 -94 68839
rect 582 68788 602 69812
rect 666 68788 686 69812
rect 582 68492 686 68788
rect -607 68440 315 68441
rect -607 67520 -606 68440
rect 314 67520 315 68440
rect -607 67519 315 67520
rect -198 67121 -94 67519
rect 582 67468 602 68492
rect 666 67468 686 68492
rect 582 67172 686 67468
rect -607 67120 315 67121
rect -607 66200 -606 67120
rect 314 66200 315 67120
rect -607 66199 315 66200
rect -198 65801 -94 66199
rect 582 66148 602 67172
rect 666 66148 686 67172
rect 582 65852 686 66148
rect -607 65800 315 65801
rect -607 64880 -606 65800
rect 314 64880 315 65800
rect -607 64879 315 64880
rect -198 64481 -94 64879
rect 582 64828 602 65852
rect 666 64828 686 65852
rect 582 64532 686 64828
rect -607 64480 315 64481
rect -607 63560 -606 64480
rect 314 63560 315 64480
rect -607 63559 315 63560
rect -198 63161 -94 63559
rect 582 63508 602 64532
rect 666 63508 686 64532
rect 582 63212 686 63508
rect -607 63160 315 63161
rect -607 62240 -606 63160
rect 314 62240 315 63160
rect -607 62239 315 62240
rect -198 61841 -94 62239
rect 582 62188 602 63212
rect 666 62188 686 63212
rect 582 61892 686 62188
rect -607 61840 315 61841
rect -607 60920 -606 61840
rect 314 60920 315 61840
rect -607 60919 315 60920
rect -198 60521 -94 60919
rect 582 60868 602 61892
rect 666 60868 686 61892
rect 582 60572 686 60868
rect -607 60520 315 60521
rect -607 59600 -606 60520
rect 314 59600 315 60520
rect -607 59599 315 59600
rect -198 59201 -94 59599
rect 582 59548 602 60572
rect 666 59548 686 60572
rect 582 59252 686 59548
rect -607 59200 315 59201
rect -607 58280 -606 59200
rect 314 58280 315 59200
rect -607 58279 315 58280
rect -198 57881 -94 58279
rect 582 58228 602 59252
rect 666 58228 686 59252
rect 582 57932 686 58228
rect -607 57880 315 57881
rect -607 56960 -606 57880
rect 314 56960 315 57880
rect -607 56959 315 56960
rect -198 56561 -94 56959
rect 582 56908 602 57932
rect 666 56908 686 57932
rect 582 56612 686 56908
rect -607 56560 315 56561
rect -607 55640 -606 56560
rect 314 55640 315 56560
rect -607 55639 315 55640
rect -198 55241 -94 55639
rect 582 55588 602 56612
rect 666 55588 686 56612
rect 582 55292 686 55588
rect -607 55240 315 55241
rect -607 54320 -606 55240
rect 314 54320 315 55240
rect -607 54319 315 54320
rect -198 53921 -94 54319
rect 582 54268 602 55292
rect 666 54268 686 55292
rect 582 53972 686 54268
rect -607 53920 315 53921
rect -607 53000 -606 53920
rect 314 53000 315 53920
rect -607 52999 315 53000
rect -198 52601 -94 52999
rect 582 52948 602 53972
rect 666 52948 686 53972
rect 582 52652 686 52948
rect -607 52600 315 52601
rect -607 51680 -606 52600
rect 314 51680 315 52600
rect -607 51679 315 51680
rect -198 51281 -94 51679
rect 582 51628 602 52652
rect 666 51628 686 52652
rect 582 51332 686 51628
rect -607 51280 315 51281
rect -607 50360 -606 51280
rect 314 50360 315 51280
rect -607 50359 315 50360
rect -198 49961 -94 50359
rect 582 50308 602 51332
rect 666 50308 686 51332
rect 582 50012 686 50308
rect -607 49960 315 49961
rect -607 49040 -606 49960
rect 314 49040 315 49960
rect -607 49039 315 49040
rect -198 48641 -94 49039
rect 582 48988 602 50012
rect 666 48988 686 50012
rect 582 48692 686 48988
rect -607 48640 315 48641
rect -607 47720 -606 48640
rect 314 47720 315 48640
rect -607 47719 315 47720
rect -198 47321 -94 47719
rect 582 47668 602 48692
rect 666 47668 686 48692
rect 582 47372 686 47668
rect -607 47320 315 47321
rect -607 46400 -606 47320
rect 314 46400 315 47320
rect -607 46399 315 46400
rect -198 46001 -94 46399
rect 582 46348 602 47372
rect 666 46348 686 47372
rect 582 46052 686 46348
rect -607 46000 315 46001
rect -607 45080 -606 46000
rect 314 45080 315 46000
rect -607 45079 315 45080
rect -198 44681 -94 45079
rect 582 45028 602 46052
rect 666 45028 686 46052
rect 582 44732 686 45028
rect -607 44680 315 44681
rect -607 43760 -606 44680
rect 314 43760 315 44680
rect -607 43759 315 43760
rect -198 43361 -94 43759
rect 582 43708 602 44732
rect 666 43708 686 44732
rect 582 43412 686 43708
rect -607 43360 315 43361
rect -607 42440 -606 43360
rect 314 42440 315 43360
rect -607 42439 315 42440
rect -198 42041 -94 42439
rect 582 42388 602 43412
rect 666 42388 686 43412
rect 582 42092 686 42388
rect -607 42040 315 42041
rect -607 41120 -606 42040
rect 314 41120 315 42040
rect -607 41119 315 41120
rect -198 40721 -94 41119
rect 582 41068 602 42092
rect 666 41068 686 42092
rect 582 40772 686 41068
rect -607 40720 315 40721
rect -607 39800 -606 40720
rect 314 39800 315 40720
rect -607 39799 315 39800
rect -198 39401 -94 39799
rect 582 39748 602 40772
rect 666 39748 686 40772
rect 582 39452 686 39748
rect -607 39400 315 39401
rect -607 38480 -606 39400
rect 314 38480 315 39400
rect -607 38479 315 38480
rect -198 38081 -94 38479
rect 582 38428 602 39452
rect 666 38428 686 39452
rect 582 38132 686 38428
rect -607 38080 315 38081
rect -607 37160 -606 38080
rect 314 37160 315 38080
rect -607 37159 315 37160
rect -198 36761 -94 37159
rect 582 37108 602 38132
rect 666 37108 686 38132
rect 582 36812 686 37108
rect -607 36760 315 36761
rect -607 35840 -606 36760
rect 314 35840 315 36760
rect -607 35839 315 35840
rect -198 35441 -94 35839
rect 582 35788 602 36812
rect 666 35788 686 36812
rect 582 35492 686 35788
rect -607 35440 315 35441
rect -607 34520 -606 35440
rect 314 34520 315 35440
rect -607 34519 315 34520
rect -198 34121 -94 34519
rect 582 34468 602 35492
rect 666 34468 686 35492
rect 582 34172 686 34468
rect -607 34120 315 34121
rect -607 33200 -606 34120
rect 314 33200 315 34120
rect -607 33199 315 33200
rect -198 32801 -94 33199
rect 582 33148 602 34172
rect 666 33148 686 34172
rect 582 32852 686 33148
rect -607 32800 315 32801
rect -607 31880 -606 32800
rect 314 31880 315 32800
rect -607 31879 315 31880
rect -198 31481 -94 31879
rect 582 31828 602 32852
rect 666 31828 686 32852
rect 582 31532 686 31828
rect -607 31480 315 31481
rect -607 30560 -606 31480
rect 314 30560 315 31480
rect -607 30559 315 30560
rect -198 30161 -94 30559
rect 582 30508 602 31532
rect 666 30508 686 31532
rect 582 30212 686 30508
rect -607 30160 315 30161
rect -607 29240 -606 30160
rect 314 29240 315 30160
rect -607 29239 315 29240
rect -198 28841 -94 29239
rect 582 29188 602 30212
rect 666 29188 686 30212
rect 582 28892 686 29188
rect -607 28840 315 28841
rect -607 27920 -606 28840
rect 314 27920 315 28840
rect -607 27919 315 27920
rect -198 27521 -94 27919
rect 582 27868 602 28892
rect 666 27868 686 28892
rect 582 27572 686 27868
rect -607 27520 315 27521
rect -607 26600 -606 27520
rect 314 26600 315 27520
rect -607 26599 315 26600
rect -198 26201 -94 26599
rect 582 26548 602 27572
rect 666 26548 686 27572
rect 582 26252 686 26548
rect -607 26200 315 26201
rect -607 25280 -606 26200
rect 314 25280 315 26200
rect -607 25279 315 25280
rect -198 24881 -94 25279
rect 582 25228 602 26252
rect 666 25228 686 26252
rect 582 24932 686 25228
rect -607 24880 315 24881
rect -607 23960 -606 24880
rect 314 23960 315 24880
rect -607 23959 315 23960
rect -198 23561 -94 23959
rect 582 23908 602 24932
rect 666 23908 686 24932
rect 582 23612 686 23908
rect -607 23560 315 23561
rect -607 22640 -606 23560
rect 314 22640 315 23560
rect -607 22639 315 22640
rect -198 22241 -94 22639
rect 582 22588 602 23612
rect 666 22588 686 23612
rect 582 22292 686 22588
rect -607 22240 315 22241
rect -607 21320 -606 22240
rect 314 21320 315 22240
rect -607 21319 315 21320
rect -198 20921 -94 21319
rect 582 21268 602 22292
rect 666 21268 686 22292
rect 582 20972 686 21268
rect -607 20920 315 20921
rect -607 20000 -606 20920
rect 314 20000 315 20920
rect -607 19999 315 20000
rect -198 19601 -94 19999
rect 582 19948 602 20972
rect 666 19948 686 20972
rect 582 19652 686 19948
rect -607 19600 315 19601
rect -607 18680 -606 19600
rect 314 18680 315 19600
rect -607 18679 315 18680
rect -198 18281 -94 18679
rect 582 18628 602 19652
rect 666 18628 686 19652
rect 582 18332 686 18628
rect -607 18280 315 18281
rect -607 17360 -606 18280
rect 314 17360 315 18280
rect -607 17359 315 17360
rect -198 16961 -94 17359
rect 582 17308 602 18332
rect 666 17308 686 18332
rect 582 17012 686 17308
rect -607 16960 315 16961
rect -607 16040 -606 16960
rect 314 16040 315 16960
rect -607 16039 315 16040
rect -198 15641 -94 16039
rect 582 15988 602 17012
rect 666 15988 686 17012
rect 582 15692 686 15988
rect -607 15640 315 15641
rect -607 14720 -606 15640
rect 314 14720 315 15640
rect -607 14719 315 14720
rect -198 14321 -94 14719
rect 582 14668 602 15692
rect 666 14668 686 15692
rect 582 14372 686 14668
rect -607 14320 315 14321
rect -607 13400 -606 14320
rect 314 13400 315 14320
rect -607 13399 315 13400
rect -198 13001 -94 13399
rect 582 13348 602 14372
rect 666 13348 686 14372
rect 582 13052 686 13348
rect -607 13000 315 13001
rect -607 12080 -606 13000
rect 314 12080 315 13000
rect -607 12079 315 12080
rect -198 11681 -94 12079
rect 582 12028 602 13052
rect 666 12028 686 13052
rect 582 11732 686 12028
rect -607 11680 315 11681
rect -607 10760 -606 11680
rect 314 10760 315 11680
rect -607 10759 315 10760
rect -198 10361 -94 10759
rect 582 10708 602 11732
rect 666 10708 686 11732
rect 582 10412 686 10708
rect -607 10360 315 10361
rect -607 9440 -606 10360
rect 314 9440 315 10360
rect -607 9439 315 9440
rect -198 9041 -94 9439
rect 582 9388 602 10412
rect 666 9388 686 10412
rect 582 9092 686 9388
rect -607 9040 315 9041
rect -607 8120 -606 9040
rect 314 8120 315 9040
rect -607 8119 315 8120
rect -198 7721 -94 8119
rect 582 8068 602 9092
rect 666 8068 686 9092
rect 582 7772 686 8068
rect -607 7720 315 7721
rect -607 6800 -606 7720
rect 314 6800 315 7720
rect -607 6799 315 6800
rect -198 6401 -94 6799
rect 582 6748 602 7772
rect 666 6748 686 7772
rect 582 6452 686 6748
rect -607 6400 315 6401
rect -607 5480 -606 6400
rect 314 5480 315 6400
rect -607 5479 315 5480
rect -198 5081 -94 5479
rect 582 5428 602 6452
rect 666 5428 686 6452
rect 582 5132 686 5428
rect -607 5080 315 5081
rect -607 4160 -606 5080
rect 314 4160 315 5080
rect -607 4159 315 4160
rect -198 3761 -94 4159
rect 582 4108 602 5132
rect 666 4108 686 5132
rect 582 3812 686 4108
rect -607 3760 315 3761
rect -607 2840 -606 3760
rect 314 2840 315 3760
rect -607 2839 315 2840
rect -198 2441 -94 2839
rect 582 2788 602 3812
rect 666 2788 686 3812
rect 582 2492 686 2788
rect -607 2440 315 2441
rect -607 1520 -606 2440
rect 314 1520 315 2440
rect -607 1519 315 1520
rect -198 1121 -94 1519
rect 582 1468 602 2492
rect 666 1468 686 2492
rect 582 1172 686 1468
rect -607 1120 315 1121
rect -607 200 -606 1120
rect 314 200 315 1120
rect -607 199 315 200
rect -198 -199 -94 199
rect 582 148 602 1172
rect 666 148 686 1172
rect 582 -148 686 148
rect -607 -200 315 -199
rect -607 -1120 -606 -200
rect 314 -1120 315 -200
rect -607 -1121 315 -1120
rect -198 -1519 -94 -1121
rect 582 -1172 602 -148
rect 666 -1172 686 -148
rect 582 -1468 686 -1172
rect -607 -1520 315 -1519
rect -607 -2440 -606 -1520
rect 314 -2440 315 -1520
rect -607 -2441 315 -2440
rect -198 -2839 -94 -2441
rect 582 -2492 602 -1468
rect 666 -2492 686 -1468
rect 582 -2788 686 -2492
rect -607 -2840 315 -2839
rect -607 -3760 -606 -2840
rect 314 -3760 315 -2840
rect -607 -3761 315 -3760
rect -198 -4159 -94 -3761
rect 582 -3812 602 -2788
rect 666 -3812 686 -2788
rect 582 -4108 686 -3812
rect -607 -4160 315 -4159
rect -607 -5080 -606 -4160
rect 314 -5080 315 -4160
rect -607 -5081 315 -5080
rect -198 -5479 -94 -5081
rect 582 -5132 602 -4108
rect 666 -5132 686 -4108
rect 582 -5428 686 -5132
rect -607 -5480 315 -5479
rect -607 -6400 -606 -5480
rect 314 -6400 315 -5480
rect -607 -6401 315 -6400
rect -198 -6799 -94 -6401
rect 582 -6452 602 -5428
rect 666 -6452 686 -5428
rect 582 -6748 686 -6452
rect -607 -6800 315 -6799
rect -607 -7720 -606 -6800
rect 314 -7720 315 -6800
rect -607 -7721 315 -7720
rect -198 -8119 -94 -7721
rect 582 -7772 602 -6748
rect 666 -7772 686 -6748
rect 582 -8068 686 -7772
rect -607 -8120 315 -8119
rect -607 -9040 -606 -8120
rect 314 -9040 315 -8120
rect -607 -9041 315 -9040
rect -198 -9439 -94 -9041
rect 582 -9092 602 -8068
rect 666 -9092 686 -8068
rect 582 -9388 686 -9092
rect -607 -9440 315 -9439
rect -607 -10360 -606 -9440
rect 314 -10360 315 -9440
rect -607 -10361 315 -10360
rect -198 -10759 -94 -10361
rect 582 -10412 602 -9388
rect 666 -10412 686 -9388
rect 582 -10708 686 -10412
rect -607 -10760 315 -10759
rect -607 -11680 -606 -10760
rect 314 -11680 315 -10760
rect -607 -11681 315 -11680
rect -198 -12079 -94 -11681
rect 582 -11732 602 -10708
rect 666 -11732 686 -10708
rect 582 -12028 686 -11732
rect -607 -12080 315 -12079
rect -607 -13000 -606 -12080
rect 314 -13000 315 -12080
rect -607 -13001 315 -13000
rect -198 -13399 -94 -13001
rect 582 -13052 602 -12028
rect 666 -13052 686 -12028
rect 582 -13348 686 -13052
rect -607 -13400 315 -13399
rect -607 -14320 -606 -13400
rect 314 -14320 315 -13400
rect -607 -14321 315 -14320
rect -198 -14719 -94 -14321
rect 582 -14372 602 -13348
rect 666 -14372 686 -13348
rect 582 -14668 686 -14372
rect -607 -14720 315 -14719
rect -607 -15640 -606 -14720
rect 314 -15640 315 -14720
rect -607 -15641 315 -15640
rect -198 -16039 -94 -15641
rect 582 -15692 602 -14668
rect 666 -15692 686 -14668
rect 582 -15988 686 -15692
rect -607 -16040 315 -16039
rect -607 -16960 -606 -16040
rect 314 -16960 315 -16040
rect -607 -16961 315 -16960
rect -198 -17359 -94 -16961
rect 582 -17012 602 -15988
rect 666 -17012 686 -15988
rect 582 -17308 686 -17012
rect -607 -17360 315 -17359
rect -607 -18280 -606 -17360
rect 314 -18280 315 -17360
rect -607 -18281 315 -18280
rect -198 -18679 -94 -18281
rect 582 -18332 602 -17308
rect 666 -18332 686 -17308
rect 582 -18628 686 -18332
rect -607 -18680 315 -18679
rect -607 -19600 -606 -18680
rect 314 -19600 315 -18680
rect -607 -19601 315 -19600
rect -198 -19999 -94 -19601
rect 582 -19652 602 -18628
rect 666 -19652 686 -18628
rect 582 -19948 686 -19652
rect -607 -20000 315 -19999
rect -607 -20920 -606 -20000
rect 314 -20920 315 -20000
rect -607 -20921 315 -20920
rect -198 -21319 -94 -20921
rect 582 -20972 602 -19948
rect 666 -20972 686 -19948
rect 582 -21268 686 -20972
rect -607 -21320 315 -21319
rect -607 -22240 -606 -21320
rect 314 -22240 315 -21320
rect -607 -22241 315 -22240
rect -198 -22639 -94 -22241
rect 582 -22292 602 -21268
rect 666 -22292 686 -21268
rect 582 -22588 686 -22292
rect -607 -22640 315 -22639
rect -607 -23560 -606 -22640
rect 314 -23560 315 -22640
rect -607 -23561 315 -23560
rect -198 -23959 -94 -23561
rect 582 -23612 602 -22588
rect 666 -23612 686 -22588
rect 582 -23908 686 -23612
rect -607 -23960 315 -23959
rect -607 -24880 -606 -23960
rect 314 -24880 315 -23960
rect -607 -24881 315 -24880
rect -198 -25279 -94 -24881
rect 582 -24932 602 -23908
rect 666 -24932 686 -23908
rect 582 -25228 686 -24932
rect -607 -25280 315 -25279
rect -607 -26200 -606 -25280
rect 314 -26200 315 -25280
rect -607 -26201 315 -26200
rect -198 -26599 -94 -26201
rect 582 -26252 602 -25228
rect 666 -26252 686 -25228
rect 582 -26548 686 -26252
rect -607 -26600 315 -26599
rect -607 -27520 -606 -26600
rect 314 -27520 315 -26600
rect -607 -27521 315 -27520
rect -198 -27919 -94 -27521
rect 582 -27572 602 -26548
rect 666 -27572 686 -26548
rect 582 -27868 686 -27572
rect -607 -27920 315 -27919
rect -607 -28840 -606 -27920
rect 314 -28840 315 -27920
rect -607 -28841 315 -28840
rect -198 -29239 -94 -28841
rect 582 -28892 602 -27868
rect 666 -28892 686 -27868
rect 582 -29188 686 -28892
rect -607 -29240 315 -29239
rect -607 -30160 -606 -29240
rect 314 -30160 315 -29240
rect -607 -30161 315 -30160
rect -198 -30559 -94 -30161
rect 582 -30212 602 -29188
rect 666 -30212 686 -29188
rect 582 -30508 686 -30212
rect -607 -30560 315 -30559
rect -607 -31480 -606 -30560
rect 314 -31480 315 -30560
rect -607 -31481 315 -31480
rect -198 -31879 -94 -31481
rect 582 -31532 602 -30508
rect 666 -31532 686 -30508
rect 582 -31828 686 -31532
rect -607 -31880 315 -31879
rect -607 -32800 -606 -31880
rect 314 -32800 315 -31880
rect -607 -32801 315 -32800
rect -198 -33199 -94 -32801
rect 582 -32852 602 -31828
rect 666 -32852 686 -31828
rect 582 -33148 686 -32852
rect -607 -33200 315 -33199
rect -607 -34120 -606 -33200
rect 314 -34120 315 -33200
rect -607 -34121 315 -34120
rect -198 -34519 -94 -34121
rect 582 -34172 602 -33148
rect 666 -34172 686 -33148
rect 582 -34468 686 -34172
rect -607 -34520 315 -34519
rect -607 -35440 -606 -34520
rect 314 -35440 315 -34520
rect -607 -35441 315 -35440
rect -198 -35839 -94 -35441
rect 582 -35492 602 -34468
rect 666 -35492 686 -34468
rect 582 -35788 686 -35492
rect -607 -35840 315 -35839
rect -607 -36760 -606 -35840
rect 314 -36760 315 -35840
rect -607 -36761 315 -36760
rect -198 -37159 -94 -36761
rect 582 -36812 602 -35788
rect 666 -36812 686 -35788
rect 582 -37108 686 -36812
rect -607 -37160 315 -37159
rect -607 -38080 -606 -37160
rect 314 -38080 315 -37160
rect -607 -38081 315 -38080
rect -198 -38479 -94 -38081
rect 582 -38132 602 -37108
rect 666 -38132 686 -37108
rect 582 -38428 686 -38132
rect -607 -38480 315 -38479
rect -607 -39400 -606 -38480
rect 314 -39400 315 -38480
rect -607 -39401 315 -39400
rect -198 -39799 -94 -39401
rect 582 -39452 602 -38428
rect 666 -39452 686 -38428
rect 582 -39748 686 -39452
rect -607 -39800 315 -39799
rect -607 -40720 -606 -39800
rect 314 -40720 315 -39800
rect -607 -40721 315 -40720
rect -198 -41119 -94 -40721
rect 582 -40772 602 -39748
rect 666 -40772 686 -39748
rect 582 -41068 686 -40772
rect -607 -41120 315 -41119
rect -607 -42040 -606 -41120
rect 314 -42040 315 -41120
rect -607 -42041 315 -42040
rect -198 -42439 -94 -42041
rect 582 -42092 602 -41068
rect 666 -42092 686 -41068
rect 582 -42388 686 -42092
rect -607 -42440 315 -42439
rect -607 -43360 -606 -42440
rect 314 -43360 315 -42440
rect -607 -43361 315 -43360
rect -198 -43759 -94 -43361
rect 582 -43412 602 -42388
rect 666 -43412 686 -42388
rect 582 -43708 686 -43412
rect -607 -43760 315 -43759
rect -607 -44680 -606 -43760
rect 314 -44680 315 -43760
rect -607 -44681 315 -44680
rect -198 -45079 -94 -44681
rect 582 -44732 602 -43708
rect 666 -44732 686 -43708
rect 582 -45028 686 -44732
rect -607 -45080 315 -45079
rect -607 -46000 -606 -45080
rect 314 -46000 315 -45080
rect -607 -46001 315 -46000
rect -198 -46399 -94 -46001
rect 582 -46052 602 -45028
rect 666 -46052 686 -45028
rect 582 -46348 686 -46052
rect -607 -46400 315 -46399
rect -607 -47320 -606 -46400
rect 314 -47320 315 -46400
rect -607 -47321 315 -47320
rect -198 -47719 -94 -47321
rect 582 -47372 602 -46348
rect 666 -47372 686 -46348
rect 582 -47668 686 -47372
rect -607 -47720 315 -47719
rect -607 -48640 -606 -47720
rect 314 -48640 315 -47720
rect -607 -48641 315 -48640
rect -198 -49039 -94 -48641
rect 582 -48692 602 -47668
rect 666 -48692 686 -47668
rect 582 -48988 686 -48692
rect -607 -49040 315 -49039
rect -607 -49960 -606 -49040
rect 314 -49960 315 -49040
rect -607 -49961 315 -49960
rect -198 -50359 -94 -49961
rect 582 -50012 602 -48988
rect 666 -50012 686 -48988
rect 582 -50308 686 -50012
rect -607 -50360 315 -50359
rect -607 -51280 -606 -50360
rect 314 -51280 315 -50360
rect -607 -51281 315 -51280
rect -198 -51679 -94 -51281
rect 582 -51332 602 -50308
rect 666 -51332 686 -50308
rect 582 -51628 686 -51332
rect -607 -51680 315 -51679
rect -607 -52600 -606 -51680
rect 314 -52600 315 -51680
rect -607 -52601 315 -52600
rect -198 -52999 -94 -52601
rect 582 -52652 602 -51628
rect 666 -52652 686 -51628
rect 582 -52948 686 -52652
rect -607 -53000 315 -52999
rect -607 -53920 -606 -53000
rect 314 -53920 315 -53000
rect -607 -53921 315 -53920
rect -198 -54319 -94 -53921
rect 582 -53972 602 -52948
rect 666 -53972 686 -52948
rect 582 -54268 686 -53972
rect -607 -54320 315 -54319
rect -607 -55240 -606 -54320
rect 314 -55240 315 -54320
rect -607 -55241 315 -55240
rect -198 -55639 -94 -55241
rect 582 -55292 602 -54268
rect 666 -55292 686 -54268
rect 582 -55588 686 -55292
rect -607 -55640 315 -55639
rect -607 -56560 -606 -55640
rect 314 -56560 315 -55640
rect -607 -56561 315 -56560
rect -198 -56959 -94 -56561
rect 582 -56612 602 -55588
rect 666 -56612 686 -55588
rect 582 -56908 686 -56612
rect -607 -56960 315 -56959
rect -607 -57880 -606 -56960
rect 314 -57880 315 -56960
rect -607 -57881 315 -57880
rect -198 -58279 -94 -57881
rect 582 -57932 602 -56908
rect 666 -57932 686 -56908
rect 582 -58228 686 -57932
rect -607 -58280 315 -58279
rect -607 -59200 -606 -58280
rect 314 -59200 315 -58280
rect -607 -59201 315 -59200
rect -198 -59599 -94 -59201
rect 582 -59252 602 -58228
rect 666 -59252 686 -58228
rect 582 -59548 686 -59252
rect -607 -59600 315 -59599
rect -607 -60520 -606 -59600
rect 314 -60520 315 -59600
rect -607 -60521 315 -60520
rect -198 -60919 -94 -60521
rect 582 -60572 602 -59548
rect 666 -60572 686 -59548
rect 582 -60868 686 -60572
rect -607 -60920 315 -60919
rect -607 -61840 -606 -60920
rect 314 -61840 315 -60920
rect -607 -61841 315 -61840
rect -198 -62239 -94 -61841
rect 582 -61892 602 -60868
rect 666 -61892 686 -60868
rect 582 -62188 686 -61892
rect -607 -62240 315 -62239
rect -607 -63160 -606 -62240
rect 314 -63160 315 -62240
rect -607 -63161 315 -63160
rect -198 -63559 -94 -63161
rect 582 -63212 602 -62188
rect 666 -63212 686 -62188
rect 582 -63508 686 -63212
rect -607 -63560 315 -63559
rect -607 -64480 -606 -63560
rect 314 -64480 315 -63560
rect -607 -64481 315 -64480
rect -198 -64879 -94 -64481
rect 582 -64532 602 -63508
rect 666 -64532 686 -63508
rect 582 -64828 686 -64532
rect -607 -64880 315 -64879
rect -607 -65800 -606 -64880
rect 314 -65800 315 -64880
rect -607 -65801 315 -65800
rect -198 -66199 -94 -65801
rect 582 -65852 602 -64828
rect 666 -65852 686 -64828
rect 582 -66148 686 -65852
rect -607 -66200 315 -66199
rect -607 -67120 -606 -66200
rect 314 -67120 315 -66200
rect -607 -67121 315 -67120
rect -198 -67519 -94 -67121
rect 582 -67172 602 -66148
rect 666 -67172 686 -66148
rect 582 -67468 686 -67172
rect -607 -67520 315 -67519
rect -607 -68440 -606 -67520
rect 314 -68440 315 -67520
rect -607 -68441 315 -68440
rect -198 -68839 -94 -68441
rect 582 -68492 602 -67468
rect 666 -68492 686 -67468
rect 582 -68788 686 -68492
rect -607 -68840 315 -68839
rect -607 -69760 -606 -68840
rect 314 -69760 315 -68840
rect -607 -69761 315 -69760
rect -198 -70159 -94 -69761
rect 582 -69812 602 -68788
rect 666 -69812 686 -68788
rect 582 -70108 686 -69812
rect -607 -70160 315 -70159
rect -607 -71080 -606 -70160
rect 314 -71080 315 -70160
rect -607 -71081 315 -71080
rect -198 -71479 -94 -71081
rect 582 -71132 602 -70108
rect 666 -71132 686 -70108
rect 582 -71428 686 -71132
rect -607 -71480 315 -71479
rect -607 -72400 -606 -71480
rect 314 -72400 315 -71480
rect -607 -72401 315 -72400
rect -198 -72799 -94 -72401
rect 582 -72452 602 -71428
rect 666 -72452 686 -71428
rect 582 -72748 686 -72452
rect -607 -72800 315 -72799
rect -607 -73720 -606 -72800
rect 314 -73720 315 -72800
rect -607 -73721 315 -73720
rect -198 -74119 -94 -73721
rect 582 -73772 602 -72748
rect 666 -73772 686 -72748
rect 582 -74068 686 -73772
rect -607 -74120 315 -74119
rect -607 -75040 -606 -74120
rect 314 -75040 315 -74120
rect -607 -75041 315 -75040
rect -198 -75439 -94 -75041
rect 582 -75092 602 -74068
rect 666 -75092 686 -74068
rect 582 -75388 686 -75092
rect -607 -75440 315 -75439
rect -607 -76360 -606 -75440
rect 314 -76360 315 -75440
rect -607 -76361 315 -76360
rect -198 -76759 -94 -76361
rect 582 -76412 602 -75388
rect 666 -76412 686 -75388
rect 582 -76708 686 -76412
rect -607 -76760 315 -76759
rect -607 -77680 -606 -76760
rect 314 -77680 315 -76760
rect -607 -77681 315 -77680
rect -198 -78079 -94 -77681
rect 582 -77732 602 -76708
rect 666 -77732 686 -76708
rect 582 -78028 686 -77732
rect -607 -78080 315 -78079
rect -607 -79000 -606 -78080
rect 314 -79000 315 -78080
rect -607 -79001 315 -79000
rect -198 -79399 -94 -79001
rect 582 -79052 602 -78028
rect 666 -79052 686 -78028
rect 582 -79348 686 -79052
rect -607 -79400 315 -79399
rect -607 -80320 -606 -79400
rect 314 -80320 315 -79400
rect -607 -80321 315 -80320
rect -198 -80719 -94 -80321
rect 582 -80372 602 -79348
rect 666 -80372 686 -79348
rect 582 -80668 686 -80372
rect -607 -80720 315 -80719
rect -607 -81640 -606 -80720
rect 314 -81640 315 -80720
rect -607 -81641 315 -81640
rect -198 -82039 -94 -81641
rect 582 -81692 602 -80668
rect 666 -81692 686 -80668
rect 582 -81988 686 -81692
rect -607 -82040 315 -82039
rect -607 -82960 -606 -82040
rect 314 -82960 315 -82040
rect -607 -82961 315 -82960
rect -198 -83359 -94 -82961
rect 582 -83012 602 -81988
rect 666 -83012 686 -81988
rect 582 -83308 686 -83012
rect -607 -83360 315 -83359
rect -607 -84280 -606 -83360
rect 314 -84280 315 -83360
rect -607 -84281 315 -84280
rect -198 -84480 -94 -84281
rect 582 -84332 602 -83308
rect 666 -84332 686 -83308
rect 582 -84480 686 -84332
<< properties >>
string FIXED_BBOX -686 83280 394 84360
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5.0 l 5.0 val 53.8 carea 2.00 cperi 0.19 nx 1 ny 128 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

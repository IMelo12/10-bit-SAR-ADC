** sch_path: /home/ttuser/Documents/SARADC/xschem/cap2/cap2.sch
**.subckt cap2 bottom top
*.ipin bottom
*.ipin top
XC12 top bottom sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=2 m=2
**.ends
.end

magic
tech sky130A
magscale 1 2
timestamp 1753737846
<< viali >>
rect 1593 21641 1627 21675
rect 3985 21641 4019 21675
rect 6561 21641 6595 21675
rect 7297 21641 7331 21675
rect 9137 21641 9171 21675
rect 11713 21641 11747 21675
rect 14289 21641 14323 21675
rect 15209 21641 15243 21675
rect 16865 21641 16899 21675
rect 17601 21641 17635 21675
rect 19441 21641 19475 21675
rect 20085 21641 20119 21675
rect 1961 21573 1995 21607
rect 4537 21573 4571 21607
rect 9689 21573 9723 21607
rect 12265 21573 12299 21607
rect 1501 21505 1535 21539
rect 2329 21505 2363 21539
rect 3893 21505 3927 21539
rect 4905 21505 4939 21539
rect 6469 21505 6503 21539
rect 7205 21505 7239 21539
rect 9045 21505 9079 21539
rect 10057 21505 10091 21539
rect 11621 21505 11655 21539
rect 12633 21505 12667 21539
rect 14197 21505 14231 21539
rect 14933 21505 14967 21539
rect 16773 21505 16807 21539
rect 17509 21505 17543 21539
rect 19349 21505 19383 21539
rect 19993 21505 20027 21539
rect 1501 21097 1535 21131
rect 12587 21097 12621 21131
rect 18843 21097 18877 21131
rect 20177 21097 20211 21131
rect 7021 20961 7055 20995
rect 10655 20961 10689 20995
rect 11161 20961 11195 20995
rect 16911 20961 16945 20995
rect 17417 20961 17451 20995
rect 1685 20893 1719 20927
rect 4445 20893 4479 20927
rect 4813 20893 4847 20927
rect 7297 20893 7331 20927
rect 7665 20893 7699 20927
rect 9654 20893 9688 20927
rect 10552 20893 10586 20927
rect 10793 20893 10827 20927
rect 14105 20893 14139 20927
rect 16808 20893 16842 20927
rect 17049 20893 17083 20927
rect 19625 20893 19659 20927
rect 3985 20825 4019 20859
rect 7849 20825 7883 20859
rect 9321 20825 9355 20859
rect 13645 20825 13679 20859
rect 13829 20825 13863 20859
rect 14381 20825 14415 20859
rect 20269 20825 20303 20859
rect 4629 20757 4663 20791
rect 5549 20757 5583 20791
rect 9045 20757 9079 20791
rect 9551 20757 9585 20791
rect 15853 20757 15887 20791
rect 19809 20757 19843 20791
rect 11023 20553 11057 20587
rect 14841 20553 14875 20587
rect 20361 20553 20395 20587
rect 18475 20485 18509 20519
rect 18889 20485 18923 20519
rect 9597 20417 9631 20451
rect 18372 20417 18406 20451
rect 3617 20349 3651 20383
rect 3893 20349 3927 20383
rect 7389 20349 7423 20383
rect 7665 20349 7699 20383
rect 9229 20349 9263 20383
rect 13093 20349 13127 20383
rect 13369 20349 13403 20383
rect 18613 20349 18647 20383
rect 5365 20213 5399 20247
rect 9137 20213 9171 20247
rect 4077 20009 4111 20043
rect 6653 20009 6687 20043
rect 8999 20009 9033 20043
rect 13921 20009 13955 20043
rect 17371 20009 17405 20043
rect 8125 19873 8159 19907
rect 15439 19873 15473 19907
rect 15945 19873 15979 19907
rect 3893 19805 3927 19839
rect 8401 19805 8435 19839
rect 9102 19805 9136 19839
rect 12173 19805 12207 19839
rect 15336 19805 15370 19839
rect 15577 19805 15611 19839
rect 18128 19805 18162 19839
rect 20361 19805 20395 19839
rect 12449 19737 12483 19771
rect 18199 19669 18233 19703
rect 20177 19669 20211 19703
rect 1409 19465 1443 19499
rect 3525 19465 3559 19499
rect 13277 19465 13311 19499
rect 19717 19465 19751 19499
rect 4997 19397 5031 19431
rect 18245 19397 18279 19431
rect 3157 19329 3191 19363
rect 8217 19329 8251 19363
rect 11529 19329 11563 19363
rect 17969 19329 18003 19363
rect 2881 19261 2915 19295
rect 5273 19261 5307 19295
rect 8493 19261 8527 19295
rect 11805 19261 11839 19295
rect 9965 19125 9999 19159
rect 2007 18921 2041 18955
rect 12081 18921 12115 18955
rect 10333 18785 10367 18819
rect 1936 18717 1970 18751
rect 5181 18717 5215 18751
rect 16532 18717 16566 18751
rect 16635 18717 16669 18751
rect 17417 18717 17451 18751
rect 17601 18717 17635 18751
rect 17785 18717 17819 18751
rect 20085 18717 20119 18751
rect 5457 18649 5491 18683
rect 10609 18649 10643 18683
rect 6929 18581 6963 18615
rect 20269 18581 20303 18615
rect 5825 18377 5859 18411
rect 8769 18377 8803 18411
rect 11069 18377 11103 18411
rect 16037 18377 16071 18411
rect 4353 18309 4387 18343
rect 9597 18309 9631 18343
rect 18153 18309 18187 18343
rect 14381 18241 14415 18275
rect 14984 18241 15018 18275
rect 15393 18241 15427 18275
rect 17877 18241 17911 18275
rect 4077 18173 4111 18207
rect 7021 18173 7055 18207
rect 7297 18173 7331 18207
rect 9321 18173 9355 18207
rect 15071 18173 15105 18207
rect 15209 18173 15243 18207
rect 15853 18173 15887 18207
rect 14565 18105 14599 18139
rect 15669 18105 15703 18139
rect 15577 18037 15611 18071
rect 19625 18037 19659 18071
rect 3295 17833 3329 17867
rect 7849 17833 7883 17867
rect 15853 17833 15887 17867
rect 19625 17833 19659 17867
rect 19855 17833 19889 17867
rect 6377 17697 6411 17731
rect 11529 17697 11563 17731
rect 13645 17697 13679 17731
rect 13921 17697 13955 17731
rect 14381 17697 14415 17731
rect 1501 17629 1535 17663
rect 1869 17629 1903 17663
rect 3617 17629 3651 17663
rect 6101 17629 6135 17663
rect 11253 17629 11287 17663
rect 13277 17629 13311 17663
rect 13553 17629 13587 17663
rect 14105 17629 14139 17663
rect 18280 17629 18314 17663
rect 18383 17629 18417 17663
rect 19257 17629 19291 17663
rect 19441 17629 19475 17663
rect 19752 17629 19786 17663
rect 20085 17629 20119 17663
rect 3433 17493 3467 17527
rect 20269 17493 20303 17527
rect 1915 17289 1949 17323
rect 10195 17289 10229 17323
rect 10701 17289 10735 17323
rect 13829 17289 13863 17323
rect 17233 17289 17267 17323
rect 18061 17289 18095 17323
rect 2018 17153 2052 17187
rect 3214 17153 3248 17187
rect 3525 17153 3559 17187
rect 8160 17153 8194 17187
rect 8263 17153 8297 17187
rect 8769 17153 8803 17187
rect 10609 17153 10643 17187
rect 11529 17153 11563 17187
rect 13645 17153 13679 17187
rect 15301 17153 15335 17187
rect 15853 17153 15887 17187
rect 16773 17153 16807 17187
rect 17417 17153 17451 17187
rect 17509 17153 17543 17187
rect 18613 17153 18647 17187
rect 8401 17085 8435 17119
rect 15393 17085 15427 17119
rect 17877 17085 17911 17119
rect 18889 17085 18923 17119
rect 11713 17017 11747 17051
rect 16037 17017 16071 17051
rect 16957 17017 16991 17051
rect 17693 17017 17727 17051
rect 3111 16949 3145 16983
rect 3341 16949 3375 16983
rect 15669 16949 15703 16983
rect 20361 16949 20395 16983
rect 8217 16745 8251 16779
rect 17141 16745 17175 16779
rect 17371 16745 17405 16779
rect 19809 16677 19843 16711
rect 2973 16609 3007 16643
rect 3341 16609 3375 16643
rect 15393 16609 15427 16643
rect 15669 16609 15703 16643
rect 3157 16541 3191 16575
rect 4296 16541 4330 16575
rect 4399 16541 4433 16575
rect 4629 16541 4663 16575
rect 4813 16541 4847 16575
rect 8033 16541 8067 16575
rect 10609 16541 10643 16575
rect 17268 16541 17302 16575
rect 20085 16473 20119 16507
rect 4997 16405 5031 16439
rect 10793 16405 10827 16439
rect 9873 16201 9907 16235
rect 20269 16201 20303 16235
rect 18797 16133 18831 16167
rect 5917 16065 5951 16099
rect 6561 16065 6595 16099
rect 9689 16065 9723 16099
rect 12173 16065 12207 16099
rect 7113 15997 7147 16031
rect 7389 15997 7423 16031
rect 8861 15997 8895 16031
rect 18521 15997 18555 16031
rect 6745 15929 6779 15963
rect 6101 15861 6135 15895
rect 12357 15861 12391 15895
rect 3203 15657 3237 15691
rect 3433 15657 3467 15691
rect 11253 15657 11287 15691
rect 13369 15657 13403 15691
rect 20085 15657 20119 15691
rect 8585 15589 8619 15623
rect 16681 15589 16715 15623
rect 1409 15521 1443 15555
rect 8953 15521 8987 15555
rect 9229 15521 9263 15555
rect 14933 15521 14967 15555
rect 15209 15521 15243 15555
rect 16773 15521 16807 15555
rect 1777 15453 1811 15487
rect 3617 15453 3651 15487
rect 3950 15453 3984 15487
rect 5089 15453 5123 15487
rect 7021 15453 7055 15487
rect 7665 15453 7699 15487
rect 8401 15453 8435 15487
rect 11069 15453 11103 15487
rect 11396 15453 11430 15487
rect 11621 15453 11655 15487
rect 13610 15453 13644 15487
rect 14172 15453 14206 15487
rect 19809 15453 19843 15487
rect 7481 15385 7515 15419
rect 11483 15385 11517 15419
rect 11897 15385 11931 15419
rect 13507 15385 13541 15419
rect 17049 15385 17083 15419
rect 19993 15385 20027 15419
rect 3847 15317 3881 15351
rect 7389 15317 7423 15351
rect 7849 15317 7883 15351
rect 10701 15317 10735 15351
rect 14243 15317 14277 15351
rect 18521 15317 18555 15351
rect 19625 15317 19659 15351
rect 1915 15113 1949 15147
rect 4859 15113 4893 15147
rect 6009 15113 6043 15147
rect 8125 15113 8159 15147
rect 8401 15113 8435 15147
rect 11897 15113 11931 15147
rect 14749 15113 14783 15147
rect 17141 15113 17175 15147
rect 18521 15113 18555 15147
rect 20361 15113 20395 15147
rect 9689 15045 9723 15079
rect 11713 15045 11747 15079
rect 13277 15045 13311 15079
rect 18889 15045 18923 15079
rect 2018 14977 2052 15011
rect 3433 14977 3467 15011
rect 6193 14977 6227 15011
rect 6377 14977 6411 15011
rect 8217 14977 8251 15011
rect 8677 14977 8711 15011
rect 12081 14977 12115 15011
rect 3065 14909 3099 14943
rect 6653 14909 6687 14943
rect 9413 14909 9447 14943
rect 11529 14909 11563 14943
rect 13001 14909 13035 14943
rect 18613 14909 18647 14943
rect 8861 14841 8895 14875
rect 18153 14841 18187 14875
rect 11161 14773 11195 14807
rect 5181 14569 5215 14603
rect 15853 14569 15887 14603
rect 17049 14569 17083 14603
rect 18061 14501 18095 14535
rect 14105 14433 14139 14467
rect 4997 14365 5031 14399
rect 14381 14297 14415 14331
rect 18429 14229 18463 14263
rect 18889 13957 18923 13991
rect 1409 13889 1443 13923
rect 2237 13889 2271 13923
rect 13312 13889 13346 13923
rect 14105 13889 14139 13923
rect 3985 13821 4019 13855
rect 7849 13821 7883 13855
rect 13415 13821 13449 13855
rect 13921 13821 13955 13855
rect 14289 13821 14323 13855
rect 18613 13821 18647 13855
rect 1593 13685 1627 13719
rect 8112 13685 8146 13719
rect 9597 13685 9631 13719
rect 20361 13685 20395 13719
rect 7849 13481 7883 13515
rect 12265 13481 12299 13515
rect 13093 13481 13127 13515
rect 17417 13481 17451 13515
rect 1685 13413 1719 13447
rect 7573 13413 7607 13447
rect 9965 13413 9999 13447
rect 20177 13413 20211 13447
rect 2237 13345 2271 13379
rect 12173 13345 12207 13379
rect 12725 13345 12759 13379
rect 14105 13345 14139 13379
rect 14381 13345 14415 13379
rect 1501 13277 1535 13311
rect 1869 13277 1903 13311
rect 4997 13277 5031 13311
rect 5457 13277 5491 13311
rect 7389 13277 7423 13311
rect 7665 13277 7699 13311
rect 9505 13277 9539 13311
rect 9781 13277 9815 13311
rect 10057 13277 10091 13311
rect 10425 13277 10459 13311
rect 12449 13277 12483 13311
rect 12541 13277 12575 13311
rect 12909 13277 12943 13311
rect 17877 13277 17911 13311
rect 20361 13277 20395 13311
rect 10701 13209 10735 13243
rect 17325 13209 17359 13243
rect 5181 13141 5215 13175
rect 5641 13141 5675 13175
rect 9689 13141 9723 13175
rect 10241 13141 10275 13175
rect 15853 13141 15887 13175
rect 18153 13141 18187 13175
rect 4905 12937 4939 12971
rect 4997 12937 5031 12971
rect 7021 12937 7055 12971
rect 11345 12937 11379 12971
rect 11989 12937 12023 12971
rect 12219 12937 12253 12971
rect 8493 12869 8527 12903
rect 4721 12801 4755 12835
rect 5181 12801 5215 12835
rect 6837 12801 6871 12835
rect 7849 12801 7883 12835
rect 10241 12801 10275 12835
rect 11161 12801 11195 12835
rect 11805 12801 11839 12835
rect 12148 12801 12182 12835
rect 16681 12801 16715 12835
rect 8217 12733 8251 12767
rect 10333 12733 10367 12767
rect 10609 12733 10643 12767
rect 16957 12733 16991 12767
rect 8033 12665 8067 12699
rect 9965 12597 9999 12631
rect 18429 12597 18463 12631
rect 4721 12393 4755 12427
rect 11970 12393 12004 12427
rect 17233 12393 17267 12427
rect 18245 12325 18279 12359
rect 11713 12257 11747 12291
rect 14381 12257 14415 12291
rect 14657 12257 14691 12291
rect 4537 12189 4571 12223
rect 4997 12189 5031 12223
rect 6377 12189 6411 12223
rect 20361 12189 20395 12223
rect 16405 12121 16439 12155
rect 4813 12053 4847 12087
rect 6193 12053 6227 12087
rect 13461 12053 13495 12087
rect 18613 12053 18647 12087
rect 20177 12053 20211 12087
rect 2605 11849 2639 11883
rect 3709 11849 3743 11883
rect 4169 11849 4203 11883
rect 12081 11849 12115 11883
rect 20361 11849 20395 11883
rect 18889 11781 18923 11815
rect 1869 11713 1903 11747
rect 2421 11713 2455 11747
rect 2881 11713 2915 11747
rect 2973 11713 3007 11747
rect 3525 11713 3559 11747
rect 3985 11713 4019 11747
rect 6009 11713 6043 11747
rect 11897 11713 11931 11747
rect 13185 11713 13219 11747
rect 1777 11645 1811 11679
rect 11713 11645 11747 11679
rect 13461 11645 13495 11679
rect 18613 11645 18647 11679
rect 2697 11577 2731 11611
rect 3157 11577 3191 11611
rect 2237 11509 2271 11543
rect 6193 11509 6227 11543
rect 14933 11509 14967 11543
rect 9597 11305 9631 11339
rect 11207 11305 11241 11339
rect 14473 11305 14507 11339
rect 9413 11237 9447 11271
rect 10425 11237 10459 11271
rect 11529 11237 11563 11271
rect 6193 11169 6227 11203
rect 6469 11169 6503 11203
rect 15393 11169 15427 11203
rect 15669 11169 15703 11203
rect 17141 11169 17175 11203
rect 2881 11101 2915 11135
rect 5917 11101 5951 11135
rect 9229 11101 9263 11135
rect 9781 11101 9815 11135
rect 9873 11101 9907 11135
rect 10241 11101 10275 11135
rect 11136 11101 11170 11135
rect 11345 11101 11379 11135
rect 14105 11101 14139 11135
rect 14289 11101 14323 11135
rect 2697 10965 2731 10999
rect 6101 10965 6135 10999
rect 7941 10965 7975 10999
rect 8677 10761 8711 10795
rect 10977 10761 11011 10795
rect 11713 10761 11747 10795
rect 13967 10761 14001 10795
rect 17141 10761 17175 10795
rect 18521 10693 18555 10727
rect 18889 10693 18923 10727
rect 2421 10625 2455 10659
rect 6377 10625 6411 10659
rect 8217 10625 8251 10659
rect 8493 10625 8527 10659
rect 11529 10625 11563 10659
rect 13896 10625 13930 10659
rect 6653 10557 6687 10591
rect 8769 10557 8803 10591
rect 9045 10557 9079 10591
rect 10793 10557 10827 10591
rect 18613 10557 18647 10591
rect 8401 10489 8435 10523
rect 10609 10489 10643 10523
rect 18153 10489 18187 10523
rect 2237 10421 2271 10455
rect 8125 10421 8159 10455
rect 10517 10421 10551 10455
rect 20361 10421 20395 10455
rect 1593 10217 1627 10251
rect 7941 10217 7975 10251
rect 9137 10217 9171 10251
rect 9919 10217 9953 10251
rect 14473 10217 14507 10251
rect 17141 10217 17175 10251
rect 4261 10149 4295 10183
rect 13185 10149 13219 10183
rect 13921 10149 13955 10183
rect 18153 10149 18187 10183
rect 20177 10149 20211 10183
rect 9413 10081 9447 10115
rect 11069 10081 11103 10115
rect 11345 10081 11379 10115
rect 11713 10081 11747 10115
rect 13277 10081 13311 10115
rect 14105 10081 14139 10115
rect 14289 10081 14323 10115
rect 14749 10081 14783 10115
rect 16497 10081 16531 10115
rect 1409 10013 1443 10047
rect 2329 10013 2363 10047
rect 4445 10013 4479 10047
rect 4686 10013 4720 10047
rect 4962 10013 4996 10047
rect 7757 10013 7791 10047
rect 9505 10013 9539 10047
rect 10022 10013 10056 10047
rect 10977 10013 11011 10047
rect 11437 10013 11471 10047
rect 13461 10013 13495 10047
rect 13553 10013 13587 10047
rect 13737 10013 13771 10047
rect 20361 10013 20395 10047
rect 1961 9945 1995 9979
rect 15025 9945 15059 9979
rect 4583 9877 4617 9911
rect 4859 9877 4893 9911
rect 18521 9877 18555 9911
rect 13323 9673 13357 9707
rect 4721 9605 4755 9639
rect 2973 9537 3007 9571
rect 12449 9537 12483 9571
rect 13220 9537 13254 9571
rect 1685 9469 1719 9503
rect 4445 9469 4479 9503
rect 6193 9469 6227 9503
rect 12633 9401 12667 9435
rect 5641 9129 5675 9163
rect 3893 8993 3927 9027
rect 4169 8993 4203 9027
rect 7113 8925 7147 8959
rect 7573 8925 7607 8959
rect 20361 8925 20395 8959
rect 6745 8857 6779 8891
rect 6653 8789 6687 8823
rect 7205 8789 7239 8823
rect 7389 8789 7423 8823
rect 20177 8789 20211 8823
rect 13369 8585 13403 8619
rect 16037 8585 16071 8619
rect 20361 8585 20395 8619
rect 18889 8517 18923 8551
rect 7297 8449 7331 8483
rect 11989 8449 12023 8483
rect 12357 8449 12391 8483
rect 13185 8449 13219 8483
rect 14105 8449 14139 8483
rect 14381 8449 14415 8483
rect 15853 8449 15887 8483
rect 16957 8449 16991 8483
rect 17233 8449 17267 8483
rect 17877 8449 17911 8483
rect 18061 8449 18095 8483
rect 18153 8449 18187 8483
rect 7757 8381 7791 8415
rect 8033 8381 8067 8415
rect 17693 8381 17727 8415
rect 18613 8381 18647 8415
rect 7481 8313 7515 8347
rect 14565 8313 14599 8347
rect 17141 8313 17175 8347
rect 9505 8245 9539 8279
rect 11805 8245 11839 8279
rect 12173 8245 12207 8279
rect 14289 8245 14323 8279
rect 17417 8245 17451 8279
rect 18337 8245 18371 8279
rect 3249 8041 3283 8075
rect 8401 8041 8435 8075
rect 11897 8041 11931 8075
rect 18061 8041 18095 8075
rect 6561 7973 6595 8007
rect 9413 7973 9447 8007
rect 9873 7973 9907 8007
rect 16221 7973 16255 8007
rect 4077 7905 4111 7939
rect 6653 7905 6687 7939
rect 6929 7905 6963 7939
rect 10149 7905 10183 7939
rect 11989 7905 12023 7939
rect 12265 7905 12299 7939
rect 14473 7905 14507 7939
rect 16313 7905 16347 7939
rect 16589 7905 16623 7939
rect 2329 7837 2363 7871
rect 2881 7837 2915 7871
rect 2973 7837 3007 7871
rect 3433 7837 3467 7871
rect 3617 7837 3651 7871
rect 3847 7837 3881 7871
rect 3950 7837 3984 7871
rect 4261 7837 4295 7871
rect 4905 7837 4939 7871
rect 5089 7837 5123 7871
rect 5227 7837 5261 7871
rect 5330 7837 5364 7871
rect 6377 7837 6411 7871
rect 8953 7837 8987 7871
rect 9229 7837 9263 7871
rect 9689 7837 9723 7871
rect 18245 7837 18279 7871
rect 4445 7769 4479 7803
rect 10425 7769 10459 7803
rect 14749 7769 14783 7803
rect 18613 7769 18647 7803
rect 2513 7701 2547 7735
rect 2697 7701 2731 7735
rect 3157 7701 3191 7735
rect 4721 7701 4755 7735
rect 9137 7701 9171 7735
rect 13737 7701 13771 7735
rect 5089 7497 5123 7531
rect 7205 7497 7239 7531
rect 10885 7497 10919 7531
rect 12449 7497 12483 7531
rect 14933 7497 14967 7531
rect 15485 7497 15519 7531
rect 16865 7497 16899 7531
rect 17693 7497 17727 7531
rect 3617 7429 3651 7463
rect 9413 7429 9447 7463
rect 11805 7429 11839 7463
rect 3249 7361 3283 7395
rect 7389 7361 7423 7395
rect 9137 7361 9171 7395
rect 11161 7361 11195 7395
rect 12265 7361 12299 7395
rect 12725 7361 12759 7395
rect 15301 7361 15335 7395
rect 16681 7361 16715 7395
rect 17325 7361 17359 7395
rect 17969 7361 18003 7395
rect 18613 7361 18647 7395
rect 2881 7293 2915 7327
rect 3341 7293 3375 7327
rect 13185 7293 13219 7327
rect 13461 7293 13495 7327
rect 17417 7293 17451 7327
rect 18889 7293 18923 7327
rect 12909 7225 12943 7259
rect 17785 7225 17819 7259
rect 1455 7157 1489 7191
rect 10977 7157 11011 7191
rect 11897 7157 11931 7191
rect 2881 6953 2915 6987
rect 2605 6817 2639 6851
rect 4629 6817 4663 6851
rect 8493 6817 8527 6851
rect 2513 6749 2547 6783
rect 6653 6749 6687 6783
rect 6745 6749 6779 6783
rect 8585 6749 8619 6783
rect 10977 6749 11011 6783
rect 14381 6749 14415 6783
rect 20361 6749 20395 6783
rect 6377 6681 6411 6715
rect 7021 6681 7055 6715
rect 8769 6613 8803 6647
rect 10793 6613 10827 6647
rect 14565 6613 14599 6647
rect 20177 6613 20211 6647
rect 6791 6409 6825 6443
rect 20361 6409 20395 6443
rect 6720 6273 6754 6307
rect 9413 6273 9447 6307
rect 17509 6273 17543 6307
rect 18613 6273 18647 6307
rect 18889 6205 18923 6239
rect 9597 6069 9631 6103
rect 17325 6069 17359 6103
rect 10977 5865 11011 5899
rect 15485 5865 15519 5899
rect 8585 5797 8619 5831
rect 15117 5797 15151 5831
rect 15761 5797 15795 5831
rect 2881 5729 2915 5763
rect 3157 5729 3191 5763
rect 9229 5729 9263 5763
rect 9505 5729 9539 5763
rect 11713 5729 11747 5763
rect 15853 5729 15887 5763
rect 18061 5729 18095 5763
rect 2789 5661 2823 5695
rect 4721 5661 4755 5695
rect 4905 5661 4939 5695
rect 5043 5661 5077 5695
rect 5146 5661 5180 5695
rect 8769 5661 8803 5695
rect 11253 5661 11287 5695
rect 11437 5661 11471 5695
rect 15577 5661 15611 5695
rect 17785 5661 17819 5695
rect 20085 5661 20119 5695
rect 16129 5593 16163 5627
rect 4537 5525 4571 5559
rect 11161 5525 11195 5559
rect 13185 5525 13219 5559
rect 14105 5525 14139 5559
rect 17601 5525 17635 5559
rect 20269 5525 20303 5559
rect 5089 5321 5123 5355
rect 5549 5321 5583 5355
rect 13645 5321 13679 5355
rect 15025 5321 15059 5355
rect 18429 5321 18463 5355
rect 3617 5253 3651 5287
rect 16313 5253 16347 5287
rect 16957 5253 16991 5287
rect 1409 5185 1443 5219
rect 5365 5185 5399 5219
rect 5825 5185 5859 5219
rect 6469 5185 6503 5219
rect 9597 5185 9631 5219
rect 18521 5185 18555 5219
rect 1777 5117 1811 5151
rect 3341 5117 3375 5151
rect 5181 5117 5215 5151
rect 5917 5117 5951 5151
rect 6745 5117 6779 5151
rect 16497 5117 16531 5151
rect 16681 5117 16715 5151
rect 18797 5117 18831 5151
rect 6193 5049 6227 5083
rect 9781 5049 9815 5083
rect 14657 5049 14691 5083
rect 3203 4981 3237 5015
rect 8217 4981 8251 5015
rect 20269 4981 20303 5015
rect 4445 4777 4479 4811
rect 5319 4777 5353 4811
rect 12265 4777 12299 4811
rect 14105 4777 14139 4811
rect 15485 4777 15519 4811
rect 3985 4709 4019 4743
rect 4813 4709 4847 4743
rect 7113 4709 7147 4743
rect 15117 4709 15151 4743
rect 4997 4641 5031 4675
rect 7757 4641 7791 4675
rect 10517 4641 10551 4675
rect 10793 4641 10827 4675
rect 3801 4573 3835 4607
rect 4261 4573 4295 4607
rect 5181 4573 5215 4607
rect 5390 4573 5424 4607
rect 6929 4573 6963 4607
rect 7481 4573 7515 4607
rect 7941 4573 7975 4607
rect 8125 4573 8159 4607
rect 8263 4573 8297 4607
rect 8366 4573 8400 4607
rect 7665 4437 7699 4471
rect 8125 4097 8159 4131
rect 8309 4097 8343 4131
rect 8518 4097 8552 4131
rect 18613 4097 18647 4131
rect 18889 4029 18923 4063
rect 7941 3961 7975 3995
rect 8447 3893 8481 3927
rect 20361 3893 20395 3927
rect 7849 3689 7883 3723
rect 20269 3621 20303 3655
rect 2881 3553 2915 3587
rect 5273 3553 5307 3587
rect 8217 3553 8251 3587
rect 10701 3553 10735 3587
rect 11069 3553 11103 3587
rect 15485 3553 15519 3587
rect 15853 3553 15887 3587
rect 3157 3485 3191 3519
rect 4997 3485 5031 3519
rect 8033 3485 8067 3519
rect 9965 3485 9999 3519
rect 10517 3485 10551 3519
rect 20085 3485 20119 3519
rect 1409 3349 1443 3383
rect 6745 3349 6779 3383
rect 9781 3349 9815 3383
rect 10241 3349 10275 3383
rect 12495 3349 12529 3383
rect 17279 3349 17313 3383
rect 13829 3145 13863 3179
rect 1685 3009 1719 3043
rect 4675 3009 4709 3043
rect 4813 3009 4847 3043
rect 6653 3009 6687 3043
rect 9321 3009 9355 3043
rect 17049 3009 17083 3043
rect 20361 3009 20395 3043
rect 2881 2941 2915 2975
rect 3249 2941 3283 2975
rect 6929 2941 6963 2975
rect 9689 2941 9723 2975
rect 12081 2941 12115 2975
rect 12357 2941 12391 2975
rect 17417 2941 17451 2975
rect 1501 2805 1535 2839
rect 4997 2805 5031 2839
rect 8401 2805 8435 2839
rect 11115 2805 11149 2839
rect 18843 2805 18877 2839
rect 20177 2805 20211 2839
rect 10747 2601 10781 2635
rect 11069 2533 11103 2567
rect 4077 2465 4111 2499
rect 5825 2465 5859 2499
rect 8953 2465 8987 2499
rect 9321 2465 9355 2499
rect 1501 2397 1535 2431
rect 1961 2397 1995 2431
rect 3249 2397 3283 2431
rect 5917 2397 5951 2431
rect 7113 2397 7147 2431
rect 8401 2397 8435 2431
rect 11253 2397 11287 2431
rect 12541 2397 12575 2431
rect 13553 2397 13587 2431
rect 15117 2397 15151 2431
rect 16129 2397 16163 2431
rect 17417 2397 17451 2431
rect 18981 2397 19015 2431
rect 19533 2397 19567 2431
rect 20269 2397 20303 2431
rect 4353 2329 4387 2363
rect 1593 2261 1627 2295
rect 2145 2261 2179 2295
rect 3433 2261 3467 2295
rect 6101 2261 6135 2295
rect 7297 2261 7331 2295
rect 8585 2261 8619 2295
rect 12357 2261 12391 2295
rect 13737 2261 13771 2295
rect 14933 2261 14967 2295
rect 16313 2261 16347 2295
rect 17601 2261 17635 2295
rect 18797 2261 18831 2295
rect 19717 2261 19751 2295
rect 20177 2261 20211 2295
<< metal1 >>
rect 1104 21786 20859 21808
rect 1104 21734 5848 21786
rect 5900 21734 5912 21786
rect 5964 21734 5976 21786
rect 6028 21734 6040 21786
rect 6092 21734 6104 21786
rect 6156 21734 10747 21786
rect 10799 21734 10811 21786
rect 10863 21734 10875 21786
rect 10927 21734 10939 21786
rect 10991 21734 11003 21786
rect 11055 21734 15646 21786
rect 15698 21734 15710 21786
rect 15762 21734 15774 21786
rect 15826 21734 15838 21786
rect 15890 21734 15902 21786
rect 15954 21734 20545 21786
rect 20597 21734 20609 21786
rect 20661 21734 20673 21786
rect 20725 21734 20737 21786
rect 20789 21734 20801 21786
rect 20853 21734 20859 21786
rect 1104 21712 20859 21734
rect 566 21632 572 21684
rect 624 21672 630 21684
rect 1581 21675 1639 21681
rect 1581 21672 1593 21675
rect 624 21644 1593 21672
rect 624 21632 630 21644
rect 1581 21641 1593 21644
rect 1627 21641 1639 21675
rect 1581 21635 1639 21641
rect 3142 21632 3148 21684
rect 3200 21672 3206 21684
rect 3973 21675 4031 21681
rect 3973 21672 3985 21675
rect 3200 21644 3985 21672
rect 3200 21632 3206 21644
rect 3973 21641 3985 21644
rect 4019 21641 4031 21675
rect 3973 21635 4031 21641
rect 5718 21632 5724 21684
rect 5776 21672 5782 21684
rect 6549 21675 6607 21681
rect 6549 21672 6561 21675
rect 5776 21644 6561 21672
rect 5776 21632 5782 21644
rect 6549 21641 6561 21644
rect 6595 21641 6607 21675
rect 6549 21635 6607 21641
rect 7006 21632 7012 21684
rect 7064 21672 7070 21684
rect 7285 21675 7343 21681
rect 7285 21672 7297 21675
rect 7064 21644 7297 21672
rect 7064 21632 7070 21644
rect 7285 21641 7297 21644
rect 7331 21641 7343 21675
rect 7285 21635 7343 21641
rect 8294 21632 8300 21684
rect 8352 21672 8358 21684
rect 9125 21675 9183 21681
rect 9125 21672 9137 21675
rect 8352 21644 9137 21672
rect 8352 21632 8358 21644
rect 9125 21641 9137 21644
rect 9171 21641 9183 21675
rect 9125 21635 9183 21641
rect 10594 21632 10600 21684
rect 10652 21672 10658 21684
rect 11701 21675 11759 21681
rect 11701 21672 11713 21675
rect 10652 21644 11713 21672
rect 10652 21632 10658 21644
rect 11701 21641 11713 21644
rect 11747 21641 11759 21675
rect 11701 21635 11759 21641
rect 13446 21632 13452 21684
rect 13504 21672 13510 21684
rect 14277 21675 14335 21681
rect 14277 21672 14289 21675
rect 13504 21644 14289 21672
rect 13504 21632 13510 21644
rect 14277 21641 14289 21644
rect 14323 21641 14335 21675
rect 14277 21635 14335 21641
rect 14734 21632 14740 21684
rect 14792 21672 14798 21684
rect 15197 21675 15255 21681
rect 15197 21672 15209 21675
rect 14792 21644 15209 21672
rect 14792 21632 14798 21644
rect 15197 21641 15209 21644
rect 15243 21641 15255 21675
rect 15197 21635 15255 21641
rect 16022 21632 16028 21684
rect 16080 21672 16086 21684
rect 16853 21675 16911 21681
rect 16853 21672 16865 21675
rect 16080 21644 16865 21672
rect 16080 21632 16086 21644
rect 16853 21641 16865 21644
rect 16899 21641 16911 21675
rect 16853 21635 16911 21641
rect 17586 21632 17592 21684
rect 17644 21632 17650 21684
rect 18598 21632 18604 21684
rect 18656 21672 18662 21684
rect 19429 21675 19487 21681
rect 19429 21672 19441 21675
rect 18656 21644 19441 21672
rect 18656 21632 18662 21644
rect 19429 21641 19441 21644
rect 19475 21641 19487 21675
rect 19429 21635 19487 21641
rect 20070 21632 20076 21684
rect 20128 21632 20134 21684
rect 1946 21564 1952 21616
rect 2004 21564 2010 21616
rect 4522 21564 4528 21616
rect 4580 21564 4586 21616
rect 9582 21564 9588 21616
rect 9640 21604 9646 21616
rect 9677 21607 9735 21613
rect 9677 21604 9689 21607
rect 9640 21576 9689 21604
rect 9640 21564 9646 21576
rect 9677 21573 9689 21576
rect 9723 21573 9735 21607
rect 9677 21567 9735 21573
rect 12158 21564 12164 21616
rect 12216 21604 12222 21616
rect 12253 21607 12311 21613
rect 12253 21604 12265 21607
rect 12216 21576 12265 21604
rect 12216 21564 12222 21576
rect 12253 21573 12265 21576
rect 12299 21573 12311 21607
rect 12253 21567 12311 21573
rect 1486 21496 1492 21548
rect 1544 21496 1550 21548
rect 2317 21539 2375 21545
rect 2317 21505 2329 21539
rect 2363 21536 2375 21539
rect 3050 21536 3056 21548
rect 2363 21508 3056 21536
rect 2363 21505 2375 21508
rect 2317 21499 2375 21505
rect 3050 21496 3056 21508
rect 3108 21496 3114 21548
rect 3786 21496 3792 21548
rect 3844 21536 3850 21548
rect 3881 21539 3939 21545
rect 3881 21536 3893 21539
rect 3844 21508 3893 21536
rect 3844 21496 3850 21508
rect 3881 21505 3893 21508
rect 3927 21505 3939 21539
rect 3881 21499 3939 21505
rect 4890 21496 4896 21548
rect 4948 21496 4954 21548
rect 5626 21496 5632 21548
rect 5684 21536 5690 21548
rect 6457 21539 6515 21545
rect 6457 21536 6469 21539
rect 5684 21508 6469 21536
rect 5684 21496 5690 21508
rect 6457 21505 6469 21508
rect 6503 21505 6515 21539
rect 6457 21499 6515 21505
rect 7190 21496 7196 21548
rect 7248 21496 7254 21548
rect 8846 21496 8852 21548
rect 8904 21536 8910 21548
rect 9033 21539 9091 21545
rect 9033 21536 9045 21539
rect 8904 21508 9045 21536
rect 8904 21496 8910 21508
rect 9033 21505 9045 21508
rect 9079 21505 9091 21539
rect 9033 21499 9091 21505
rect 10042 21496 10048 21548
rect 10100 21496 10106 21548
rect 11606 21496 11612 21548
rect 11664 21496 11670 21548
rect 12618 21496 12624 21548
rect 12676 21496 12682 21548
rect 14182 21496 14188 21548
rect 14240 21496 14246 21548
rect 14921 21539 14979 21545
rect 14921 21505 14933 21539
rect 14967 21536 14979 21539
rect 15010 21536 15016 21548
rect 14967 21508 15016 21536
rect 14967 21505 14979 21508
rect 14921 21499 14979 21505
rect 15010 21496 15016 21508
rect 15068 21496 15074 21548
rect 16758 21496 16764 21548
rect 16816 21496 16822 21548
rect 17494 21496 17500 21548
rect 17552 21496 17558 21548
rect 19334 21496 19340 21548
rect 19392 21496 19398 21548
rect 19702 21496 19708 21548
rect 19760 21536 19766 21548
rect 19981 21539 20039 21545
rect 19981 21536 19993 21539
rect 19760 21508 19993 21536
rect 19760 21496 19766 21508
rect 19981 21505 19993 21508
rect 20027 21505 20039 21539
rect 19981 21499 20039 21505
rect 1104 21242 20700 21264
rect 1104 21190 3399 21242
rect 3451 21190 3463 21242
rect 3515 21190 3527 21242
rect 3579 21190 3591 21242
rect 3643 21190 3655 21242
rect 3707 21190 8298 21242
rect 8350 21190 8362 21242
rect 8414 21190 8426 21242
rect 8478 21190 8490 21242
rect 8542 21190 8554 21242
rect 8606 21190 13197 21242
rect 13249 21190 13261 21242
rect 13313 21190 13325 21242
rect 13377 21190 13389 21242
rect 13441 21190 13453 21242
rect 13505 21190 18096 21242
rect 18148 21190 18160 21242
rect 18212 21190 18224 21242
rect 18276 21190 18288 21242
rect 18340 21190 18352 21242
rect 18404 21190 20700 21242
rect 1104 21168 20700 21190
rect 1302 21088 1308 21140
rect 1360 21128 1366 21140
rect 12618 21137 12624 21140
rect 1489 21131 1547 21137
rect 1489 21128 1501 21131
rect 1360 21100 1501 21128
rect 1360 21088 1366 21100
rect 1489 21097 1501 21100
rect 1535 21097 1547 21131
rect 12575 21131 12624 21137
rect 1489 21091 1547 21097
rect 10520 21100 12480 21128
rect 7009 20995 7067 21001
rect 7009 20961 7021 20995
rect 7055 20992 7067 20995
rect 8938 20992 8944 21004
rect 7055 20964 8944 20992
rect 7055 20961 7067 20964
rect 7009 20955 7067 20961
rect 8938 20952 8944 20964
rect 8996 20952 9002 21004
rect 1673 20927 1731 20933
rect 1673 20893 1685 20927
rect 1719 20924 1731 20927
rect 4433 20927 4491 20933
rect 1719 20896 2774 20924
rect 1719 20893 1731 20896
rect 1673 20887 1731 20893
rect 2746 20856 2774 20896
rect 4433 20893 4445 20927
rect 4479 20924 4491 20927
rect 4479 20896 4660 20924
rect 4479 20893 4491 20896
rect 4433 20887 4491 20893
rect 3970 20856 3976 20868
rect 2746 20828 3976 20856
rect 3970 20816 3976 20828
rect 4028 20816 4034 20868
rect 4632 20797 4660 20896
rect 4798 20884 4804 20936
rect 4856 20884 4862 20936
rect 7282 20884 7288 20936
rect 7340 20924 7346 20936
rect 7653 20927 7711 20933
rect 7653 20924 7665 20927
rect 7340 20896 7665 20924
rect 7340 20884 7346 20896
rect 7653 20893 7665 20896
rect 7699 20924 7711 20927
rect 8202 20924 8208 20936
rect 7699 20896 8208 20924
rect 7699 20893 7711 20896
rect 7653 20887 7711 20893
rect 8202 20884 8208 20896
rect 8260 20884 8266 20936
rect 9642 20927 9700 20933
rect 9642 20893 9654 20927
rect 9688 20924 9700 20927
rect 9766 20924 9772 20936
rect 9688 20896 9772 20924
rect 9688 20893 9700 20896
rect 9642 20887 9700 20893
rect 9766 20884 9772 20896
rect 9824 20884 9830 20936
rect 10520 20933 10548 21100
rect 10643 20995 10701 21001
rect 10643 20961 10655 20995
rect 10689 20992 10701 20995
rect 11149 20995 11207 21001
rect 11149 20992 11161 20995
rect 10689 20964 11161 20992
rect 10689 20961 10701 20964
rect 10643 20955 10701 20961
rect 11149 20961 11161 20964
rect 11195 20961 11207 20995
rect 12452 20992 12480 21100
rect 12575 21097 12587 21131
rect 12621 21097 12624 21131
rect 12575 21091 12624 21097
rect 12618 21088 12624 21091
rect 12676 21088 12682 21140
rect 18831 21131 18889 21137
rect 18831 21097 18843 21131
rect 18877 21128 18889 21131
rect 19334 21128 19340 21140
rect 18877 21100 19340 21128
rect 18877 21097 18889 21100
rect 18831 21091 18889 21097
rect 19334 21088 19340 21100
rect 19392 21088 19398 21140
rect 20165 21131 20223 21137
rect 20165 21097 20177 21131
rect 20211 21128 20223 21131
rect 21174 21128 21180 21140
rect 20211 21100 21180 21128
rect 20211 21097 20223 21100
rect 20165 21091 20223 21097
rect 21174 21088 21180 21100
rect 21232 21088 21238 21140
rect 15378 20992 15384 21004
rect 12452 20964 15384 20992
rect 11149 20955 11207 20961
rect 15378 20952 15384 20964
rect 15436 20992 15442 21004
rect 16899 20995 16957 21001
rect 15436 20964 16574 20992
rect 15436 20952 15442 20964
rect 10520 20927 10598 20933
rect 10520 20896 10552 20927
rect 10540 20893 10552 20896
rect 10586 20893 10598 20927
rect 10540 20887 10598 20893
rect 10781 20927 10839 20933
rect 10781 20893 10793 20927
rect 10827 20893 10839 20927
rect 14093 20927 14151 20933
rect 14093 20924 14105 20927
rect 10781 20887 10839 20893
rect 13648 20896 14105 20924
rect 6730 20856 6736 20868
rect 6578 20828 6736 20856
rect 6730 20816 6736 20828
rect 6788 20816 6794 20868
rect 7834 20816 7840 20868
rect 7892 20816 7898 20868
rect 9306 20816 9312 20868
rect 9364 20816 9370 20868
rect 4617 20791 4675 20797
rect 4617 20757 4629 20791
rect 4663 20757 4675 20791
rect 4617 20751 4675 20757
rect 5074 20748 5080 20800
rect 5132 20788 5138 20800
rect 5537 20791 5595 20797
rect 5537 20788 5549 20791
rect 5132 20760 5549 20788
rect 5132 20748 5138 20760
rect 5537 20757 5549 20760
rect 5583 20757 5595 20791
rect 5537 20751 5595 20757
rect 9030 20748 9036 20800
rect 9088 20748 9094 20800
rect 9582 20797 9588 20800
rect 9539 20791 9588 20797
rect 9539 20757 9551 20791
rect 9585 20757 9588 20791
rect 9539 20751 9588 20757
rect 9582 20748 9588 20751
rect 9640 20748 9646 20800
rect 10502 20748 10508 20800
rect 10560 20788 10566 20800
rect 10796 20788 10824 20887
rect 12526 20856 12532 20868
rect 12190 20828 12532 20856
rect 12526 20816 12532 20828
rect 12584 20816 12590 20868
rect 13078 20816 13084 20868
rect 13136 20856 13142 20868
rect 13648 20865 13676 20896
rect 14093 20893 14105 20896
rect 14139 20893 14151 20927
rect 16546 20924 16574 20964
rect 16899 20961 16911 20995
rect 16945 20992 16957 20995
rect 17405 20995 17463 21001
rect 17405 20992 17417 20995
rect 16945 20964 17417 20992
rect 16945 20961 16957 20964
rect 16899 20955 16957 20961
rect 17405 20961 17417 20964
rect 17451 20961 17463 20995
rect 17405 20955 17463 20961
rect 16796 20927 16854 20933
rect 16796 20924 16808 20927
rect 16546 20896 16808 20924
rect 14093 20887 14151 20893
rect 16796 20893 16808 20896
rect 16842 20893 16854 20927
rect 16796 20887 16854 20893
rect 17034 20884 17040 20936
rect 17092 20884 17098 20936
rect 19610 20884 19616 20936
rect 19668 20884 19674 20936
rect 13633 20859 13691 20865
rect 13633 20856 13645 20859
rect 13136 20828 13645 20856
rect 13136 20816 13142 20828
rect 13633 20825 13645 20828
rect 13679 20825 13691 20859
rect 13633 20819 13691 20825
rect 13814 20816 13820 20868
rect 13872 20816 13878 20868
rect 14366 20816 14372 20868
rect 14424 20816 14430 20868
rect 18966 20856 18972 20868
rect 15594 20828 16574 20856
rect 18446 20828 18972 20856
rect 10560 20760 10824 20788
rect 10560 20748 10566 20760
rect 15194 20748 15200 20800
rect 15252 20788 15258 20800
rect 15841 20791 15899 20797
rect 15841 20788 15853 20791
rect 15252 20760 15853 20788
rect 15252 20748 15258 20760
rect 15841 20757 15853 20760
rect 15887 20757 15899 20791
rect 16546 20788 16574 20828
rect 18966 20816 18972 20828
rect 19024 20816 19030 20868
rect 20162 20856 20168 20868
rect 19076 20828 20168 20856
rect 19076 20788 19104 20828
rect 20162 20816 20168 20828
rect 20220 20816 20226 20868
rect 20254 20816 20260 20868
rect 20312 20816 20318 20868
rect 16546 20760 19104 20788
rect 15841 20751 15899 20757
rect 19426 20748 19432 20800
rect 19484 20788 19490 20800
rect 19797 20791 19855 20797
rect 19797 20788 19809 20791
rect 19484 20760 19809 20788
rect 19484 20748 19490 20760
rect 19797 20757 19809 20760
rect 19843 20757 19855 20791
rect 19797 20751 19855 20757
rect 1104 20698 20859 20720
rect 1104 20646 5848 20698
rect 5900 20646 5912 20698
rect 5964 20646 5976 20698
rect 6028 20646 6040 20698
rect 6092 20646 6104 20698
rect 6156 20646 10747 20698
rect 10799 20646 10811 20698
rect 10863 20646 10875 20698
rect 10927 20646 10939 20698
rect 10991 20646 11003 20698
rect 11055 20646 15646 20698
rect 15698 20646 15710 20698
rect 15762 20646 15774 20698
rect 15826 20646 15838 20698
rect 15890 20646 15902 20698
rect 15954 20646 20545 20698
rect 20597 20646 20609 20698
rect 20661 20646 20673 20698
rect 20725 20646 20737 20698
rect 20789 20646 20801 20698
rect 20853 20646 20859 20698
rect 1104 20624 20859 20646
rect 11011 20587 11069 20593
rect 11011 20553 11023 20587
rect 11057 20584 11069 20587
rect 11606 20584 11612 20596
rect 11057 20556 11612 20584
rect 11057 20553 11069 20556
rect 11011 20547 11069 20553
rect 11606 20544 11612 20556
rect 11664 20544 11670 20596
rect 14366 20544 14372 20596
rect 14424 20584 14430 20596
rect 14829 20587 14887 20593
rect 14829 20584 14841 20587
rect 14424 20556 14841 20584
rect 14424 20544 14430 20556
rect 14829 20553 14841 20556
rect 14875 20553 14887 20587
rect 14829 20547 14887 20553
rect 20254 20544 20260 20596
rect 20312 20584 20318 20596
rect 20349 20587 20407 20593
rect 20349 20584 20361 20587
rect 20312 20556 20361 20584
rect 20312 20544 20318 20556
rect 20349 20553 20361 20556
rect 20395 20553 20407 20587
rect 20349 20547 20407 20553
rect 6730 20516 6736 20528
rect 5106 20488 6736 20516
rect 6730 20476 6736 20488
rect 6788 20476 6794 20528
rect 9030 20516 9036 20528
rect 8878 20488 9036 20516
rect 9030 20476 9036 20488
rect 9088 20476 9094 20528
rect 9950 20476 9956 20528
rect 10008 20476 10014 20528
rect 12802 20476 12808 20528
rect 12860 20516 12866 20528
rect 18463 20519 18521 20525
rect 12860 20488 13846 20516
rect 12860 20476 12866 20488
rect 18463 20485 18475 20519
rect 18509 20516 18521 20519
rect 18877 20519 18935 20525
rect 18877 20516 18889 20519
rect 18509 20488 18889 20516
rect 18509 20485 18521 20488
rect 18463 20479 18521 20485
rect 18877 20485 18889 20488
rect 18923 20485 18935 20519
rect 18877 20479 18935 20485
rect 19610 20476 19616 20528
rect 19668 20476 19674 20528
rect 9582 20408 9588 20460
rect 9640 20408 9646 20460
rect 18322 20408 18328 20460
rect 18380 20457 18386 20460
rect 18380 20451 18418 20457
rect 18406 20417 18418 20451
rect 18380 20411 18418 20417
rect 18380 20408 18386 20411
rect 3605 20383 3663 20389
rect 3605 20349 3617 20383
rect 3651 20380 3663 20383
rect 3881 20383 3939 20389
rect 3651 20352 3740 20380
rect 3651 20349 3663 20352
rect 3605 20343 3663 20349
rect 3712 20244 3740 20352
rect 3881 20349 3893 20383
rect 3927 20380 3939 20383
rect 4246 20380 4252 20392
rect 3927 20352 4252 20380
rect 3927 20349 3939 20352
rect 3881 20343 3939 20349
rect 4246 20340 4252 20352
rect 4304 20380 4310 20392
rect 5074 20380 5080 20392
rect 4304 20352 5080 20380
rect 4304 20340 4310 20352
rect 5074 20340 5080 20352
rect 5132 20340 5138 20392
rect 7006 20340 7012 20392
rect 7064 20380 7070 20392
rect 7282 20380 7288 20392
rect 7064 20352 7288 20380
rect 7064 20340 7070 20352
rect 7282 20340 7288 20352
rect 7340 20380 7346 20392
rect 7377 20383 7435 20389
rect 7377 20380 7389 20383
rect 7340 20352 7389 20380
rect 7340 20340 7346 20352
rect 7377 20349 7389 20352
rect 7423 20349 7435 20383
rect 7377 20343 7435 20349
rect 7650 20340 7656 20392
rect 7708 20340 7714 20392
rect 9217 20383 9275 20389
rect 9217 20349 9229 20383
rect 9263 20380 9275 20383
rect 9398 20380 9404 20392
rect 9263 20352 9404 20380
rect 9263 20349 9275 20352
rect 9217 20343 9275 20349
rect 9398 20340 9404 20352
rect 9456 20340 9462 20392
rect 11514 20340 11520 20392
rect 11572 20380 11578 20392
rect 13078 20380 13084 20392
rect 11572 20352 13084 20380
rect 11572 20340 11578 20352
rect 13078 20340 13084 20352
rect 13136 20340 13142 20392
rect 13357 20383 13415 20389
rect 13357 20349 13369 20383
rect 13403 20380 13415 20383
rect 13906 20380 13912 20392
rect 13403 20352 13912 20380
rect 13403 20349 13415 20352
rect 13357 20343 13415 20349
rect 13906 20340 13912 20352
rect 13964 20340 13970 20392
rect 17954 20340 17960 20392
rect 18012 20380 18018 20392
rect 18601 20383 18659 20389
rect 18601 20380 18613 20383
rect 18012 20352 18613 20380
rect 18012 20340 18018 20352
rect 18601 20349 18613 20352
rect 18647 20349 18659 20383
rect 18601 20343 18659 20349
rect 4062 20244 4068 20256
rect 3712 20216 4068 20244
rect 4062 20204 4068 20216
rect 4120 20204 4126 20256
rect 5350 20204 5356 20256
rect 5408 20204 5414 20256
rect 9122 20204 9128 20256
rect 9180 20204 9186 20256
rect 16482 20204 16488 20256
rect 16540 20244 16546 20256
rect 16666 20244 16672 20256
rect 16540 20216 16672 20244
rect 16540 20204 16546 20216
rect 16666 20204 16672 20216
rect 16724 20204 16730 20256
rect 1104 20154 20700 20176
rect 1104 20102 3399 20154
rect 3451 20102 3463 20154
rect 3515 20102 3527 20154
rect 3579 20102 3591 20154
rect 3643 20102 3655 20154
rect 3707 20102 8298 20154
rect 8350 20102 8362 20154
rect 8414 20102 8426 20154
rect 8478 20102 8490 20154
rect 8542 20102 8554 20154
rect 8606 20102 13197 20154
rect 13249 20102 13261 20154
rect 13313 20102 13325 20154
rect 13377 20102 13389 20154
rect 13441 20102 13453 20154
rect 13505 20102 18096 20154
rect 18148 20102 18160 20154
rect 18212 20102 18224 20154
rect 18276 20102 18288 20154
rect 18340 20102 18352 20154
rect 18404 20102 20700 20154
rect 1104 20080 20700 20102
rect 4065 20043 4123 20049
rect 4065 20009 4077 20043
rect 4111 20040 4123 20043
rect 4798 20040 4804 20052
rect 4111 20012 4804 20040
rect 4111 20009 4123 20012
rect 4065 20003 4123 20009
rect 4798 20000 4804 20012
rect 4856 20000 4862 20052
rect 6641 20043 6699 20049
rect 6641 20009 6653 20043
rect 6687 20040 6699 20043
rect 7650 20040 7656 20052
rect 6687 20012 7656 20040
rect 6687 20009 6699 20012
rect 6641 20003 6699 20009
rect 7650 20000 7656 20012
rect 7708 20000 7714 20052
rect 8938 20000 8944 20052
rect 8996 20049 9002 20052
rect 8996 20043 9045 20049
rect 8996 20009 8999 20043
rect 9033 20009 9045 20043
rect 8996 20003 9045 20009
rect 8996 20000 9002 20003
rect 13906 20000 13912 20052
rect 13964 20000 13970 20052
rect 17359 20043 17417 20049
rect 17359 20009 17371 20043
rect 17405 20040 17417 20043
rect 17494 20040 17500 20052
rect 17405 20012 17500 20040
rect 17405 20009 17417 20012
rect 17359 20003 17417 20009
rect 17494 20000 17500 20012
rect 17552 20000 17558 20052
rect 8113 19907 8171 19913
rect 8113 19873 8125 19907
rect 8159 19904 8171 19907
rect 15194 19904 15200 19916
rect 8159 19876 15200 19904
rect 8159 19873 8171 19876
rect 8113 19867 8171 19873
rect 15194 19864 15200 19876
rect 15252 19864 15258 19916
rect 15427 19907 15485 19913
rect 15427 19873 15439 19907
rect 15473 19904 15485 19907
rect 15933 19907 15991 19913
rect 15933 19904 15945 19907
rect 15473 19876 15945 19904
rect 15473 19873 15485 19876
rect 15427 19867 15485 19873
rect 15933 19873 15945 19876
rect 15979 19873 15991 19907
rect 15933 19867 15991 19873
rect 16040 19876 17816 19904
rect 3881 19839 3939 19845
rect 3881 19805 3893 19839
rect 3927 19836 3939 19839
rect 4246 19836 4252 19848
rect 3927 19808 4252 19836
rect 3927 19805 3939 19808
rect 3881 19799 3939 19805
rect 4246 19796 4252 19808
rect 4304 19796 4310 19848
rect 8386 19796 8392 19848
rect 8444 19796 8450 19848
rect 9122 19845 9128 19848
rect 9090 19839 9128 19845
rect 9090 19805 9102 19839
rect 9090 19799 9128 19805
rect 9122 19796 9128 19799
rect 9180 19796 9186 19848
rect 11514 19796 11520 19848
rect 11572 19836 11578 19848
rect 12161 19839 12219 19845
rect 12161 19836 12173 19839
rect 11572 19808 12173 19836
rect 11572 19796 11578 19808
rect 12161 19805 12173 19808
rect 12207 19805 12219 19839
rect 12161 19799 12219 19805
rect 15286 19796 15292 19848
rect 15344 19845 15350 19848
rect 15344 19839 15382 19845
rect 15370 19836 15382 19839
rect 15370 19808 15516 19836
rect 15370 19805 15382 19808
rect 15344 19799 15382 19805
rect 15344 19796 15350 19799
rect 8938 19768 8944 19780
rect 7682 19740 8944 19768
rect 8938 19728 8944 19740
rect 8996 19728 9002 19780
rect 12434 19728 12440 19780
rect 12492 19728 12498 19780
rect 15488 19768 15516 19808
rect 15562 19796 15568 19848
rect 15620 19796 15626 19848
rect 16040 19836 16068 19876
rect 15672 19808 16068 19836
rect 17788 19836 17816 19876
rect 18116 19839 18174 19845
rect 18116 19836 18128 19839
rect 17788 19808 18128 19836
rect 15672 19768 15700 19808
rect 18116 19805 18128 19808
rect 18162 19836 18174 19839
rect 18414 19836 18420 19848
rect 18162 19808 18420 19836
rect 18162 19805 18174 19808
rect 18116 19799 18174 19805
rect 18414 19796 18420 19808
rect 18472 19796 18478 19848
rect 20346 19796 20352 19848
rect 20404 19796 20410 19848
rect 12820 19740 12926 19768
rect 15488 19740 15700 19768
rect 12820 19712 12848 19740
rect 16666 19728 16672 19780
rect 16724 19728 16730 19780
rect 18064 19740 20208 19768
rect 12802 19660 12808 19712
rect 12860 19660 12866 19712
rect 13814 19660 13820 19712
rect 13872 19700 13878 19712
rect 18064 19700 18092 19740
rect 18230 19709 18236 19712
rect 13872 19672 18092 19700
rect 18187 19703 18236 19709
rect 13872 19660 13878 19672
rect 18187 19669 18199 19703
rect 18233 19669 18236 19703
rect 18187 19663 18236 19669
rect 18230 19660 18236 19663
rect 18288 19660 18294 19712
rect 20180 19709 20208 19740
rect 20165 19703 20223 19709
rect 20165 19669 20177 19703
rect 20211 19669 20223 19703
rect 20165 19663 20223 19669
rect 1104 19610 20859 19632
rect 1104 19558 5848 19610
rect 5900 19558 5912 19610
rect 5964 19558 5976 19610
rect 6028 19558 6040 19610
rect 6092 19558 6104 19610
rect 6156 19558 10747 19610
rect 10799 19558 10811 19610
rect 10863 19558 10875 19610
rect 10927 19558 10939 19610
rect 10991 19558 11003 19610
rect 11055 19558 15646 19610
rect 15698 19558 15710 19610
rect 15762 19558 15774 19610
rect 15826 19558 15838 19610
rect 15890 19558 15902 19610
rect 15954 19558 20545 19610
rect 20597 19558 20609 19610
rect 20661 19558 20673 19610
rect 20725 19558 20737 19610
rect 20789 19558 20801 19610
rect 20853 19558 20859 19610
rect 1104 19536 20859 19558
rect 1397 19499 1455 19505
rect 1397 19465 1409 19499
rect 1443 19496 1455 19499
rect 1486 19496 1492 19508
rect 1443 19468 1492 19496
rect 1443 19465 1455 19468
rect 1397 19459 1455 19465
rect 1486 19456 1492 19468
rect 1544 19456 1550 19508
rect 3513 19499 3571 19505
rect 3513 19465 3525 19499
rect 3559 19496 3571 19499
rect 4338 19496 4344 19508
rect 3559 19468 4344 19496
rect 3559 19465 3571 19468
rect 3513 19459 3571 19465
rect 4338 19456 4344 19468
rect 4396 19456 4402 19508
rect 6730 19496 6736 19508
rect 4908 19468 6736 19496
rect 2130 19388 2136 19440
rect 2188 19388 2194 19440
rect 2958 19388 2964 19440
rect 3016 19428 3022 19440
rect 4908 19428 4936 19468
rect 6730 19456 6736 19468
rect 6788 19456 6794 19508
rect 12434 19456 12440 19508
rect 12492 19496 12498 19508
rect 13265 19499 13323 19505
rect 13265 19496 13277 19499
rect 12492 19468 13277 19496
rect 12492 19456 12498 19468
rect 13265 19465 13277 19468
rect 13311 19465 13323 19499
rect 13265 19459 13323 19465
rect 19702 19456 19708 19508
rect 19760 19456 19766 19508
rect 3016 19400 3188 19428
rect 4554 19400 4936 19428
rect 4985 19431 5043 19437
rect 3016 19388 3022 19400
rect 3160 19369 3188 19400
rect 4985 19397 4997 19431
rect 5031 19428 5043 19431
rect 5350 19428 5356 19440
rect 5031 19400 5356 19428
rect 5031 19397 5043 19400
rect 4985 19391 5043 19397
rect 5350 19388 5356 19400
rect 5408 19388 5414 19440
rect 9030 19388 9036 19440
rect 9088 19388 9094 19440
rect 12802 19388 12808 19440
rect 12860 19388 12866 19440
rect 18230 19388 18236 19440
rect 18288 19388 18294 19440
rect 18782 19388 18788 19440
rect 18840 19388 18846 19440
rect 3145 19363 3203 19369
rect 3145 19329 3157 19363
rect 3191 19329 3203 19363
rect 3145 19323 3203 19329
rect 7834 19320 7840 19372
rect 7892 19360 7898 19372
rect 8018 19360 8024 19372
rect 7892 19332 8024 19360
rect 7892 19320 7898 19332
rect 8018 19320 8024 19332
rect 8076 19360 8082 19372
rect 8205 19363 8263 19369
rect 8205 19360 8217 19363
rect 8076 19332 8217 19360
rect 8076 19320 8082 19332
rect 8205 19329 8217 19332
rect 8251 19329 8263 19363
rect 8205 19323 8263 19329
rect 10318 19320 10324 19372
rect 10376 19360 10382 19372
rect 11514 19360 11520 19372
rect 10376 19332 11520 19360
rect 10376 19320 10382 19332
rect 11514 19320 11520 19332
rect 11572 19320 11578 19372
rect 17954 19320 17960 19372
rect 18012 19320 18018 19372
rect 2866 19252 2872 19304
rect 2924 19252 2930 19304
rect 5261 19295 5319 19301
rect 5261 19292 5273 19295
rect 5184 19264 5273 19292
rect 5184 19168 5212 19264
rect 5261 19261 5273 19264
rect 5307 19261 5319 19295
rect 5261 19255 5319 19261
rect 8481 19295 8539 19301
rect 8481 19261 8493 19295
rect 8527 19292 8539 19295
rect 8846 19292 8852 19304
rect 8527 19264 8852 19292
rect 8527 19261 8539 19264
rect 8481 19255 8539 19261
rect 8846 19252 8852 19264
rect 8904 19252 8910 19304
rect 11790 19252 11796 19304
rect 11848 19252 11854 19304
rect 5166 19116 5172 19168
rect 5224 19116 5230 19168
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 9953 19159 10011 19165
rect 9953 19156 9965 19159
rect 9732 19128 9965 19156
rect 9732 19116 9738 19128
rect 9953 19125 9965 19128
rect 9999 19125 10011 19159
rect 9953 19119 10011 19125
rect 1104 19066 20700 19088
rect 1104 19014 3399 19066
rect 3451 19014 3463 19066
rect 3515 19014 3527 19066
rect 3579 19014 3591 19066
rect 3643 19014 3655 19066
rect 3707 19014 8298 19066
rect 8350 19014 8362 19066
rect 8414 19014 8426 19066
rect 8478 19014 8490 19066
rect 8542 19014 8554 19066
rect 8606 19014 13197 19066
rect 13249 19014 13261 19066
rect 13313 19014 13325 19066
rect 13377 19014 13389 19066
rect 13441 19014 13453 19066
rect 13505 19014 18096 19066
rect 18148 19014 18160 19066
rect 18212 19014 18224 19066
rect 18276 19014 18288 19066
rect 18340 19014 18352 19066
rect 18404 19014 20700 19066
rect 1104 18992 20700 19014
rect 1995 18955 2053 18961
rect 1995 18921 2007 18955
rect 2041 18952 2053 18955
rect 2866 18952 2872 18964
rect 2041 18924 2872 18952
rect 2041 18921 2053 18924
rect 1995 18915 2053 18921
rect 2866 18912 2872 18924
rect 2924 18912 2930 18964
rect 11790 18912 11796 18964
rect 11848 18952 11854 18964
rect 12069 18955 12127 18961
rect 12069 18952 12081 18955
rect 11848 18924 12081 18952
rect 11848 18912 11854 18924
rect 12069 18921 12081 18924
rect 12115 18921 12127 18955
rect 12069 18915 12127 18921
rect 8018 18776 8024 18828
rect 8076 18816 8082 18828
rect 10318 18816 10324 18828
rect 8076 18788 10324 18816
rect 8076 18776 8082 18788
rect 10318 18776 10324 18788
rect 10376 18776 10382 18828
rect 1946 18757 1952 18760
rect 1924 18751 1952 18757
rect 1924 18717 1936 18751
rect 1924 18711 1952 18717
rect 1946 18708 1952 18711
rect 2004 18708 2010 18760
rect 4062 18708 4068 18760
rect 4120 18748 4126 18760
rect 5166 18748 5172 18760
rect 4120 18720 5172 18748
rect 4120 18708 4126 18720
rect 5166 18708 5172 18720
rect 5224 18708 5230 18760
rect 16022 18708 16028 18760
rect 16080 18748 16086 18760
rect 16520 18751 16578 18757
rect 16520 18748 16532 18751
rect 16080 18720 16532 18748
rect 16080 18708 16086 18720
rect 16520 18717 16532 18720
rect 16566 18717 16578 18751
rect 16520 18711 16578 18717
rect 16623 18751 16681 18757
rect 16623 18717 16635 18751
rect 16669 18748 16681 18751
rect 17405 18751 17463 18757
rect 17405 18748 17417 18751
rect 16669 18720 17417 18748
rect 16669 18717 16681 18720
rect 16623 18711 16681 18717
rect 17405 18717 17417 18720
rect 17451 18717 17463 18751
rect 17405 18711 17463 18717
rect 17586 18708 17592 18760
rect 17644 18708 17650 18760
rect 17773 18751 17831 18757
rect 17773 18717 17785 18751
rect 17819 18748 17831 18751
rect 18782 18748 18788 18760
rect 17819 18720 18788 18748
rect 17819 18717 17831 18720
rect 17773 18711 17831 18717
rect 18782 18708 18788 18720
rect 18840 18708 18846 18760
rect 20070 18708 20076 18760
rect 20128 18708 20134 18760
rect 5445 18683 5503 18689
rect 5445 18649 5457 18683
rect 5491 18680 5503 18683
rect 5718 18680 5724 18692
rect 5491 18652 5724 18680
rect 5491 18649 5503 18652
rect 5445 18643 5503 18649
rect 5718 18640 5724 18652
rect 5776 18640 5782 18692
rect 6730 18680 6736 18692
rect 6670 18652 6736 18680
rect 6730 18640 6736 18652
rect 6788 18640 6794 18692
rect 10594 18640 10600 18692
rect 10652 18640 10658 18692
rect 10704 18652 11086 18680
rect 6914 18572 6920 18624
rect 6972 18572 6978 18624
rect 9306 18572 9312 18624
rect 9364 18612 9370 18624
rect 10704 18612 10732 18652
rect 9364 18584 10732 18612
rect 10980 18612 11008 18652
rect 12802 18612 12808 18624
rect 10980 18584 12808 18612
rect 9364 18572 9370 18584
rect 12802 18572 12808 18584
rect 12860 18572 12866 18624
rect 20254 18572 20260 18624
rect 20312 18572 20318 18624
rect 1104 18522 20859 18544
rect 1104 18470 5848 18522
rect 5900 18470 5912 18522
rect 5964 18470 5976 18522
rect 6028 18470 6040 18522
rect 6092 18470 6104 18522
rect 6156 18470 10747 18522
rect 10799 18470 10811 18522
rect 10863 18470 10875 18522
rect 10927 18470 10939 18522
rect 10991 18470 11003 18522
rect 11055 18470 15646 18522
rect 15698 18470 15710 18522
rect 15762 18470 15774 18522
rect 15826 18470 15838 18522
rect 15890 18470 15902 18522
rect 15954 18470 20545 18522
rect 20597 18470 20609 18522
rect 20661 18470 20673 18522
rect 20725 18470 20737 18522
rect 20789 18470 20801 18522
rect 20853 18470 20859 18522
rect 1104 18448 20859 18470
rect 5718 18368 5724 18420
rect 5776 18408 5782 18420
rect 5813 18411 5871 18417
rect 5813 18408 5825 18411
rect 5776 18380 5825 18408
rect 5776 18368 5782 18380
rect 5813 18377 5825 18380
rect 5859 18377 5871 18411
rect 5813 18371 5871 18377
rect 8757 18411 8815 18417
rect 8757 18377 8769 18411
rect 8803 18408 8815 18411
rect 8846 18408 8852 18420
rect 8803 18380 8852 18408
rect 8803 18377 8815 18380
rect 8757 18371 8815 18377
rect 8846 18368 8852 18380
rect 8904 18368 8910 18420
rect 9306 18368 9312 18420
rect 9364 18408 9370 18420
rect 9364 18380 9812 18408
rect 9364 18368 9370 18380
rect 4338 18300 4344 18352
rect 4396 18300 4402 18352
rect 6730 18340 6736 18352
rect 5566 18312 6736 18340
rect 6730 18300 6736 18312
rect 6788 18300 6794 18352
rect 9030 18340 9036 18352
rect 8510 18312 9036 18340
rect 9030 18300 9036 18312
rect 9088 18300 9094 18352
rect 9585 18343 9643 18349
rect 9585 18309 9597 18343
rect 9631 18340 9643 18343
rect 9674 18340 9680 18352
rect 9631 18312 9680 18340
rect 9631 18309 9643 18312
rect 9585 18303 9643 18309
rect 9674 18300 9680 18312
rect 9732 18300 9738 18352
rect 9784 18340 9812 18380
rect 10594 18368 10600 18420
rect 10652 18408 10658 18420
rect 11057 18411 11115 18417
rect 11057 18408 11069 18411
rect 10652 18380 11069 18408
rect 10652 18368 10658 18380
rect 11057 18377 11069 18380
rect 11103 18377 11115 18411
rect 11057 18371 11115 18377
rect 16022 18368 16028 18420
rect 16080 18368 16086 18420
rect 15654 18340 15660 18352
rect 9784 18312 10074 18340
rect 15304 18312 15660 18340
rect 14366 18232 14372 18284
rect 14424 18232 14430 18284
rect 14972 18275 15030 18281
rect 14972 18241 14984 18275
rect 15018 18272 15030 18275
rect 15304 18272 15332 18312
rect 15654 18300 15660 18312
rect 15712 18300 15718 18352
rect 18141 18343 18199 18349
rect 18141 18309 18153 18343
rect 18187 18340 18199 18343
rect 18414 18340 18420 18352
rect 18187 18312 18420 18340
rect 18187 18309 18199 18312
rect 18141 18303 18199 18309
rect 18414 18300 18420 18312
rect 18472 18300 18478 18352
rect 18782 18300 18788 18352
rect 18840 18300 18846 18352
rect 15018 18244 15332 18272
rect 15381 18275 15439 18281
rect 15018 18241 15030 18244
rect 14972 18235 15030 18241
rect 15381 18241 15393 18275
rect 15427 18241 15439 18275
rect 15381 18235 15439 18241
rect 4062 18164 4068 18216
rect 4120 18164 4126 18216
rect 7006 18164 7012 18216
rect 7064 18164 7070 18216
rect 7285 18207 7343 18213
rect 7285 18173 7297 18207
rect 7331 18204 7343 18207
rect 7834 18204 7840 18216
rect 7331 18176 7840 18204
rect 7331 18173 7343 18176
rect 7285 18167 7343 18173
rect 7834 18164 7840 18176
rect 7892 18164 7898 18216
rect 8018 18164 8024 18216
rect 8076 18204 8082 18216
rect 9309 18207 9367 18213
rect 9309 18204 9321 18207
rect 8076 18176 9321 18204
rect 8076 18164 8082 18176
rect 9309 18173 9321 18176
rect 9355 18173 9367 18207
rect 9309 18167 9367 18173
rect 15059 18207 15117 18213
rect 15059 18173 15071 18207
rect 15105 18204 15117 18207
rect 15197 18207 15255 18213
rect 15197 18204 15209 18207
rect 15105 18176 15209 18204
rect 15105 18173 15117 18176
rect 15059 18167 15117 18173
rect 15197 18173 15209 18176
rect 15243 18173 15255 18207
rect 15197 18167 15255 18173
rect 15396 18204 15424 18235
rect 17862 18232 17868 18284
rect 17920 18232 17926 18284
rect 15841 18207 15899 18213
rect 15841 18204 15853 18207
rect 15396 18176 15853 18204
rect 14553 18139 14611 18145
rect 14553 18105 14565 18139
rect 14599 18136 14611 18139
rect 15396 18136 15424 18176
rect 15841 18173 15853 18176
rect 15887 18173 15899 18207
rect 15841 18167 15899 18173
rect 14599 18108 15424 18136
rect 14599 18105 14611 18108
rect 14553 18099 14611 18105
rect 15654 18096 15660 18148
rect 15712 18096 15718 18148
rect 15286 18028 15292 18080
rect 15344 18068 15350 18080
rect 15562 18068 15568 18080
rect 15344 18040 15568 18068
rect 15344 18028 15350 18040
rect 15562 18028 15568 18040
rect 15620 18028 15626 18080
rect 19518 18028 19524 18080
rect 19576 18068 19582 18080
rect 19613 18071 19671 18077
rect 19613 18068 19625 18071
rect 19576 18040 19625 18068
rect 19576 18028 19582 18040
rect 19613 18037 19625 18040
rect 19659 18037 19671 18071
rect 19613 18031 19671 18037
rect 1104 17978 20700 18000
rect 1104 17926 3399 17978
rect 3451 17926 3463 17978
rect 3515 17926 3527 17978
rect 3579 17926 3591 17978
rect 3643 17926 3655 17978
rect 3707 17926 8298 17978
rect 8350 17926 8362 17978
rect 8414 17926 8426 17978
rect 8478 17926 8490 17978
rect 8542 17926 8554 17978
rect 8606 17926 13197 17978
rect 13249 17926 13261 17978
rect 13313 17926 13325 17978
rect 13377 17926 13389 17978
rect 13441 17926 13453 17978
rect 13505 17926 18096 17978
rect 18148 17926 18160 17978
rect 18212 17926 18224 17978
rect 18276 17926 18288 17978
rect 18340 17926 18352 17978
rect 18404 17926 20700 17978
rect 1104 17904 20700 17926
rect 3283 17867 3341 17873
rect 3283 17833 3295 17867
rect 3329 17864 3341 17867
rect 3786 17864 3792 17876
rect 3329 17836 3792 17864
rect 3329 17833 3341 17836
rect 3283 17827 3341 17833
rect 3786 17824 3792 17836
rect 3844 17824 3850 17876
rect 7006 17864 7012 17876
rect 6104 17836 7012 17864
rect 1486 17620 1492 17672
rect 1544 17620 1550 17672
rect 1854 17620 1860 17672
rect 1912 17620 1918 17672
rect 3605 17663 3663 17669
rect 3605 17629 3617 17663
rect 3651 17660 3663 17663
rect 4062 17660 4068 17672
rect 3651 17632 4068 17660
rect 3651 17629 3663 17632
rect 3605 17623 3663 17629
rect 4062 17620 4068 17632
rect 4120 17660 4126 17672
rect 6104 17669 6132 17836
rect 7006 17824 7012 17836
rect 7064 17824 7070 17876
rect 7834 17824 7840 17876
rect 7892 17824 7898 17876
rect 9950 17824 9956 17876
rect 10008 17864 10014 17876
rect 10008 17836 15516 17864
rect 10008 17824 10014 17836
rect 6365 17731 6423 17737
rect 6365 17697 6377 17731
rect 6411 17728 6423 17731
rect 6914 17728 6920 17740
rect 6411 17700 6920 17728
rect 6411 17697 6423 17700
rect 6365 17691 6423 17697
rect 6914 17688 6920 17700
rect 6972 17688 6978 17740
rect 11517 17731 11575 17737
rect 11517 17697 11529 17731
rect 11563 17728 11575 17731
rect 13633 17731 13691 17737
rect 13633 17728 13645 17731
rect 11563 17700 13645 17728
rect 11563 17697 11575 17700
rect 11517 17691 11575 17697
rect 13633 17697 13645 17700
rect 13679 17728 13691 17731
rect 13722 17728 13728 17740
rect 13679 17700 13728 17728
rect 13679 17697 13691 17700
rect 13633 17691 13691 17697
rect 13722 17688 13728 17700
rect 13780 17688 13786 17740
rect 13909 17731 13967 17737
rect 13909 17697 13921 17731
rect 13955 17728 13967 17731
rect 14369 17731 14427 17737
rect 14369 17728 14381 17731
rect 13955 17700 14381 17728
rect 13955 17697 13967 17700
rect 13909 17691 13967 17697
rect 14369 17697 14381 17700
rect 14415 17697 14427 17731
rect 14369 17691 14427 17697
rect 6089 17663 6147 17669
rect 6089 17660 6101 17663
rect 4120 17632 6101 17660
rect 4120 17620 4126 17632
rect 6089 17629 6101 17632
rect 6135 17629 6147 17663
rect 6089 17623 6147 17629
rect 11241 17663 11299 17669
rect 11241 17629 11253 17663
rect 11287 17629 11299 17663
rect 11241 17623 11299 17629
rect 13265 17663 13323 17669
rect 13265 17629 13277 17663
rect 13311 17660 13323 17663
rect 13538 17660 13544 17672
rect 13311 17632 13544 17660
rect 13311 17629 13323 17632
rect 13265 17623 13323 17629
rect 2866 17552 2872 17604
rect 2924 17592 2930 17604
rect 9030 17592 9036 17604
rect 2924 17564 3004 17592
rect 7590 17564 9036 17592
rect 2924 17552 2930 17564
rect 2130 17484 2136 17536
rect 2188 17524 2194 17536
rect 2976 17524 3004 17564
rect 2188 17496 3004 17524
rect 3421 17527 3479 17533
rect 2188 17484 2194 17496
rect 3421 17493 3433 17527
rect 3467 17524 3479 17527
rect 3510 17524 3516 17536
rect 3467 17496 3516 17524
rect 3467 17493 3479 17496
rect 3421 17487 3479 17493
rect 3510 17484 3516 17496
rect 3568 17484 3574 17536
rect 6730 17484 6736 17536
rect 6788 17524 6794 17536
rect 7668 17524 7696 17564
rect 9030 17552 9036 17564
rect 9088 17552 9094 17604
rect 11256 17536 11284 17623
rect 13538 17620 13544 17632
rect 13596 17620 13602 17672
rect 14090 17620 14096 17672
rect 14148 17620 14154 17672
rect 15488 17660 15516 17836
rect 15654 17824 15660 17876
rect 15712 17864 15718 17876
rect 15841 17867 15899 17873
rect 15841 17864 15853 17867
rect 15712 17836 15853 17864
rect 15712 17824 15718 17836
rect 15841 17833 15853 17836
rect 15887 17833 15899 17867
rect 15841 17827 15899 17833
rect 19610 17824 19616 17876
rect 19668 17824 19674 17876
rect 19843 17867 19901 17873
rect 19843 17833 19855 17867
rect 19889 17864 19901 17867
rect 20070 17864 20076 17876
rect 19889 17836 20076 17864
rect 19889 17833 19901 17836
rect 19843 17827 19901 17833
rect 20070 17824 20076 17836
rect 20128 17824 20134 17876
rect 17586 17688 17592 17740
rect 17644 17728 17650 17740
rect 17644 17700 19472 17728
rect 17644 17688 17650 17700
rect 16482 17660 16488 17672
rect 15488 17646 16488 17660
rect 15502 17632 16488 17646
rect 16482 17620 16488 17632
rect 16540 17620 16546 17672
rect 18046 17620 18052 17672
rect 18104 17660 18110 17672
rect 19444 17669 19472 17700
rect 18268 17663 18326 17669
rect 18268 17660 18280 17663
rect 18104 17632 18280 17660
rect 18104 17620 18110 17632
rect 18268 17629 18280 17632
rect 18314 17629 18326 17663
rect 18268 17623 18326 17629
rect 18371 17663 18429 17669
rect 18371 17629 18383 17663
rect 18417 17660 18429 17663
rect 19245 17663 19303 17669
rect 19245 17660 19257 17663
rect 18417 17632 19257 17660
rect 18417 17629 18429 17632
rect 18371 17623 18429 17629
rect 19245 17629 19257 17632
rect 19291 17629 19303 17663
rect 19245 17623 19303 17629
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17629 19487 17663
rect 19740 17663 19798 17669
rect 19740 17660 19752 17663
rect 19429 17623 19487 17629
rect 19536 17632 19752 17660
rect 12526 17552 12532 17604
rect 12584 17552 12590 17604
rect 18506 17552 18512 17604
rect 18564 17592 18570 17604
rect 19536 17592 19564 17632
rect 19740 17629 19752 17632
rect 19786 17629 19798 17663
rect 19740 17623 19798 17629
rect 20070 17620 20076 17672
rect 20128 17620 20134 17672
rect 18564 17564 19564 17592
rect 18564 17552 18570 17564
rect 6788 17496 7696 17524
rect 6788 17484 6794 17496
rect 11238 17484 11244 17536
rect 11296 17524 11302 17536
rect 17954 17524 17960 17536
rect 11296 17496 17960 17524
rect 11296 17484 11302 17496
rect 17954 17484 17960 17496
rect 18012 17484 18018 17536
rect 20254 17484 20260 17536
rect 20312 17484 20318 17536
rect 1104 17434 20859 17456
rect 1104 17382 5848 17434
rect 5900 17382 5912 17434
rect 5964 17382 5976 17434
rect 6028 17382 6040 17434
rect 6092 17382 6104 17434
rect 6156 17382 10747 17434
rect 10799 17382 10811 17434
rect 10863 17382 10875 17434
rect 10927 17382 10939 17434
rect 10991 17382 11003 17434
rect 11055 17382 15646 17434
rect 15698 17382 15710 17434
rect 15762 17382 15774 17434
rect 15826 17382 15838 17434
rect 15890 17382 15902 17434
rect 15954 17382 20545 17434
rect 20597 17382 20609 17434
rect 20661 17382 20673 17434
rect 20725 17382 20737 17434
rect 20789 17382 20801 17434
rect 20853 17382 20859 17434
rect 1104 17360 20859 17382
rect 1854 17280 1860 17332
rect 1912 17329 1918 17332
rect 1912 17323 1961 17329
rect 1912 17289 1915 17323
rect 1949 17289 1961 17323
rect 1912 17283 1961 17289
rect 1912 17280 1918 17283
rect 2866 17280 2872 17332
rect 2924 17320 2930 17332
rect 2924 17292 9904 17320
rect 2924 17280 2930 17292
rect 9876 17252 9904 17292
rect 10042 17280 10048 17332
rect 10100 17320 10106 17332
rect 10183 17323 10241 17329
rect 10183 17320 10195 17323
rect 10100 17292 10195 17320
rect 10100 17280 10106 17292
rect 10183 17289 10195 17292
rect 10229 17289 10241 17323
rect 10183 17283 10241 17289
rect 10689 17323 10747 17329
rect 10689 17289 10701 17323
rect 10735 17320 10747 17323
rect 11238 17320 11244 17332
rect 10735 17292 11244 17320
rect 10735 17289 10747 17292
rect 10689 17283 10747 17289
rect 11238 17280 11244 17292
rect 11296 17280 11302 17332
rect 13817 17323 13875 17329
rect 13817 17289 13829 17323
rect 13863 17320 13875 17323
rect 14366 17320 14372 17332
rect 13863 17292 14372 17320
rect 13863 17289 13875 17292
rect 13817 17283 13875 17289
rect 14366 17280 14372 17292
rect 14424 17280 14430 17332
rect 17034 17280 17040 17332
rect 17092 17320 17098 17332
rect 17218 17320 17224 17332
rect 17092 17292 17224 17320
rect 17092 17280 17098 17292
rect 17218 17280 17224 17292
rect 17276 17280 17282 17332
rect 18046 17280 18052 17332
rect 18104 17280 18110 17332
rect 9950 17252 9956 17264
rect 9798 17224 9956 17252
rect 9950 17212 9956 17224
rect 10008 17212 10014 17264
rect 13538 17212 13544 17264
rect 13596 17252 13602 17264
rect 17678 17252 17684 17264
rect 13596 17224 17684 17252
rect 13596 17212 13602 17224
rect 1946 17144 1952 17196
rect 2004 17193 2010 17196
rect 2004 17187 2064 17193
rect 2004 17153 2018 17187
rect 2052 17184 2064 17187
rect 3202 17187 3260 17193
rect 2052 17156 2774 17184
rect 2052 17153 2064 17156
rect 2004 17147 2064 17153
rect 2004 17144 2010 17147
rect 2746 17048 2774 17156
rect 3202 17153 3214 17187
rect 3248 17184 3260 17187
rect 3248 17156 3464 17184
rect 3248 17153 3260 17156
rect 3202 17147 3260 17153
rect 3436 17116 3464 17156
rect 3510 17144 3516 17196
rect 3568 17144 3574 17196
rect 8148 17187 8206 17193
rect 8148 17184 8160 17187
rect 8128 17153 8160 17184
rect 8194 17153 8206 17187
rect 8128 17147 8206 17153
rect 8251 17187 8309 17193
rect 8251 17153 8263 17187
rect 8297 17184 8309 17187
rect 8757 17187 8815 17193
rect 8757 17184 8769 17187
rect 8297 17156 8769 17184
rect 8297 17153 8309 17156
rect 8251 17147 8309 17153
rect 8757 17153 8769 17156
rect 8803 17153 8815 17187
rect 8757 17147 8815 17153
rect 3786 17116 3792 17128
rect 3436 17088 3792 17116
rect 3786 17076 3792 17088
rect 3844 17076 3850 17128
rect 8128 17116 8156 17147
rect 9582 17144 9588 17196
rect 9640 17184 9646 17196
rect 10597 17187 10655 17193
rect 10597 17184 10609 17187
rect 9640 17156 10609 17184
rect 9640 17144 9646 17156
rect 10597 17153 10609 17156
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17153 11575 17187
rect 11517 17147 11575 17153
rect 13633 17187 13691 17193
rect 13633 17153 13645 17187
rect 13679 17184 13691 17187
rect 14090 17184 14096 17196
rect 13679 17156 14096 17184
rect 13679 17153 13691 17156
rect 13633 17147 13691 17153
rect 8389 17119 8447 17125
rect 8128 17088 8248 17116
rect 2746 17020 4016 17048
rect 3988 16992 4016 17020
rect 3142 16989 3148 16992
rect 3099 16983 3148 16989
rect 3099 16949 3111 16983
rect 3145 16949 3148 16983
rect 3099 16943 3148 16949
rect 3142 16940 3148 16943
rect 3200 16940 3206 16992
rect 3234 16940 3240 16992
rect 3292 16980 3298 16992
rect 3329 16983 3387 16989
rect 3329 16980 3341 16983
rect 3292 16952 3341 16980
rect 3292 16940 3298 16952
rect 3329 16949 3341 16952
rect 3375 16949 3387 16983
rect 3329 16943 3387 16949
rect 3970 16940 3976 16992
rect 4028 16980 4034 16992
rect 8220 16980 8248 17088
rect 8389 17085 8401 17119
rect 8435 17116 8447 17119
rect 9490 17116 9496 17128
rect 8435 17088 9496 17116
rect 8435 17085 8447 17088
rect 8389 17079 8447 17085
rect 9490 17076 9496 17088
rect 9548 17076 9554 17128
rect 9766 17076 9772 17128
rect 9824 17116 9830 17128
rect 11532 17116 11560 17147
rect 14090 17144 14096 17156
rect 14148 17184 14154 17196
rect 14918 17184 14924 17196
rect 14148 17156 14924 17184
rect 14148 17144 14154 17156
rect 14918 17144 14924 17156
rect 14976 17144 14982 17196
rect 15304 17193 15332 17224
rect 17678 17212 17684 17224
rect 17736 17212 17742 17264
rect 19610 17212 19616 17264
rect 19668 17212 19674 17264
rect 15289 17187 15347 17193
rect 15289 17153 15301 17187
rect 15335 17153 15347 17187
rect 15289 17147 15347 17153
rect 15470 17144 15476 17196
rect 15528 17184 15534 17196
rect 15841 17187 15899 17193
rect 15841 17184 15853 17187
rect 15528 17156 15853 17184
rect 15528 17144 15534 17156
rect 15841 17153 15853 17156
rect 15887 17153 15899 17187
rect 16761 17187 16819 17193
rect 16761 17184 16773 17187
rect 15841 17147 15899 17153
rect 16546 17156 16773 17184
rect 13722 17116 13728 17128
rect 9824 17088 11560 17116
rect 12406 17088 13728 17116
rect 9824 17076 9830 17088
rect 11701 17051 11759 17057
rect 11701 17017 11713 17051
rect 11747 17048 11759 17051
rect 12406 17048 12434 17088
rect 13722 17076 13728 17088
rect 13780 17116 13786 17128
rect 15381 17119 15439 17125
rect 15381 17116 15393 17119
rect 13780 17088 15393 17116
rect 13780 17076 13786 17088
rect 15381 17085 15393 17088
rect 15427 17116 15439 17119
rect 15427 17088 15792 17116
rect 15427 17085 15439 17088
rect 15381 17079 15439 17085
rect 11747 17020 12434 17048
rect 11747 17017 11759 17020
rect 11701 17011 11759 17017
rect 9766 16980 9772 16992
rect 4028 16952 9772 16980
rect 4028 16940 4034 16952
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 15654 16940 15660 16992
rect 15712 16940 15718 16992
rect 15764 16980 15792 17088
rect 16025 17051 16083 17057
rect 16025 17017 16037 17051
rect 16071 17048 16083 17051
rect 16546 17048 16574 17156
rect 16761 17153 16773 17156
rect 16807 17153 16819 17187
rect 17405 17187 17463 17193
rect 17405 17184 17417 17187
rect 16761 17147 16819 17153
rect 16960 17156 17417 17184
rect 16960 17057 16988 17156
rect 17405 17153 17417 17156
rect 17451 17153 17463 17187
rect 17405 17147 17463 17153
rect 17420 17116 17448 17147
rect 17494 17144 17500 17196
rect 17552 17144 17558 17196
rect 17954 17144 17960 17196
rect 18012 17184 18018 17196
rect 18601 17187 18659 17193
rect 18601 17184 18613 17187
rect 18012 17156 18613 17184
rect 18012 17144 18018 17156
rect 18601 17153 18613 17156
rect 18647 17153 18659 17187
rect 18601 17147 18659 17153
rect 17865 17119 17923 17125
rect 17865 17116 17877 17119
rect 17420 17088 17877 17116
rect 17865 17085 17877 17088
rect 17911 17085 17923 17119
rect 18877 17119 18935 17125
rect 18877 17116 18889 17119
rect 17865 17079 17923 17085
rect 18708 17088 18889 17116
rect 16071 17020 16574 17048
rect 16945 17051 17003 17057
rect 16071 17017 16083 17020
rect 16025 17011 16083 17017
rect 16945 17017 16957 17051
rect 16991 17017 17003 17051
rect 16945 17011 17003 17017
rect 17126 17008 17132 17060
rect 17184 17048 17190 17060
rect 17681 17051 17739 17057
rect 17681 17048 17693 17051
rect 17184 17020 17693 17048
rect 17184 17008 17190 17020
rect 17681 17017 17693 17020
rect 17727 17017 17739 17051
rect 17681 17011 17739 17017
rect 18414 16980 18420 16992
rect 15764 16952 18420 16980
rect 18414 16940 18420 16952
rect 18472 16980 18478 16992
rect 18708 16980 18736 17088
rect 18877 17085 18889 17088
rect 18923 17085 18935 17119
rect 18877 17079 18935 17085
rect 18472 16952 18736 16980
rect 20349 16983 20407 16989
rect 18472 16940 18478 16952
rect 20349 16949 20361 16983
rect 20395 16980 20407 16983
rect 20438 16980 20444 16992
rect 20395 16952 20444 16980
rect 20395 16949 20407 16952
rect 20349 16943 20407 16949
rect 20438 16940 20444 16952
rect 20496 16940 20502 16992
rect 1104 16890 20700 16912
rect 1104 16838 3399 16890
rect 3451 16838 3463 16890
rect 3515 16838 3527 16890
rect 3579 16838 3591 16890
rect 3643 16838 3655 16890
rect 3707 16838 8298 16890
rect 8350 16838 8362 16890
rect 8414 16838 8426 16890
rect 8478 16838 8490 16890
rect 8542 16838 8554 16890
rect 8606 16838 13197 16890
rect 13249 16838 13261 16890
rect 13313 16838 13325 16890
rect 13377 16838 13389 16890
rect 13441 16838 13453 16890
rect 13505 16838 18096 16890
rect 18148 16838 18160 16890
rect 18212 16838 18224 16890
rect 18276 16838 18288 16890
rect 18340 16838 18352 16890
rect 18404 16838 20700 16890
rect 1104 16816 20700 16838
rect 8205 16779 8263 16785
rect 8205 16745 8217 16779
rect 8251 16776 8263 16779
rect 9582 16776 9588 16788
rect 8251 16748 9588 16776
rect 8251 16745 8263 16748
rect 8205 16739 8263 16745
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 12802 16736 12808 16788
rect 12860 16776 12866 16788
rect 12860 16748 17080 16776
rect 12860 16736 12866 16748
rect 17052 16708 17080 16748
rect 17126 16736 17132 16788
rect 17184 16736 17190 16788
rect 17359 16779 17417 16785
rect 17359 16745 17371 16779
rect 17405 16776 17417 16779
rect 17494 16776 17500 16788
rect 17405 16748 17500 16776
rect 17405 16745 17417 16748
rect 17359 16739 17417 16745
rect 17494 16736 17500 16748
rect 17552 16736 17558 16788
rect 19797 16711 19855 16717
rect 19797 16708 19809 16711
rect 17052 16680 19809 16708
rect 19797 16677 19809 16680
rect 19843 16708 19855 16711
rect 19886 16708 19892 16720
rect 19843 16680 19892 16708
rect 19843 16677 19855 16680
rect 19797 16671 19855 16677
rect 19886 16668 19892 16680
rect 19944 16668 19950 16720
rect 2866 16600 2872 16652
rect 2924 16640 2930 16652
rect 2961 16643 3019 16649
rect 2961 16640 2973 16643
rect 2924 16612 2973 16640
rect 2924 16600 2930 16612
rect 2961 16609 2973 16612
rect 3007 16609 3019 16643
rect 2961 16603 3019 16609
rect 3234 16600 3240 16652
rect 3292 16640 3298 16652
rect 3329 16643 3387 16649
rect 3329 16640 3341 16643
rect 3292 16612 3341 16640
rect 3292 16600 3298 16612
rect 3329 16609 3341 16612
rect 3375 16609 3387 16643
rect 9306 16640 9312 16652
rect 3329 16603 3387 16609
rect 4816 16612 9312 16640
rect 3142 16532 3148 16584
rect 3200 16532 3206 16584
rect 3786 16532 3792 16584
rect 3844 16572 3850 16584
rect 4816 16581 4844 16612
rect 9306 16600 9312 16612
rect 9364 16600 9370 16652
rect 15378 16640 15384 16652
rect 15359 16612 15384 16640
rect 15378 16600 15384 16612
rect 15436 16600 15442 16652
rect 15654 16600 15660 16652
rect 15712 16600 15718 16652
rect 4284 16575 4342 16581
rect 4284 16572 4296 16575
rect 3844 16544 4296 16572
rect 3844 16532 3850 16544
rect 4284 16541 4296 16544
rect 4330 16541 4342 16575
rect 4284 16535 4342 16541
rect 4387 16575 4445 16581
rect 4387 16541 4399 16575
rect 4433 16572 4445 16575
rect 4617 16575 4675 16581
rect 4617 16572 4629 16575
rect 4433 16544 4629 16572
rect 4433 16541 4445 16544
rect 4387 16535 4445 16541
rect 4617 16541 4629 16544
rect 4663 16541 4675 16575
rect 4617 16535 4675 16541
rect 4801 16575 4859 16581
rect 4801 16541 4813 16575
rect 4847 16541 4859 16575
rect 4801 16535 4859 16541
rect 8018 16532 8024 16584
rect 8076 16532 8082 16584
rect 9858 16532 9864 16584
rect 9916 16572 9922 16584
rect 10597 16575 10655 16581
rect 10597 16572 10609 16575
rect 9916 16544 10609 16572
rect 9916 16532 9922 16544
rect 10597 16541 10609 16544
rect 10643 16541 10655 16575
rect 10597 16535 10655 16541
rect 4982 16396 4988 16448
rect 5040 16396 5046 16448
rect 10781 16439 10839 16445
rect 10781 16405 10793 16439
rect 10827 16436 10839 16439
rect 15396 16436 15424 16600
rect 10827 16408 15424 16436
rect 10827 16405 10839 16408
rect 10781 16399 10839 16405
rect 16574 16396 16580 16448
rect 16632 16436 16638 16448
rect 16776 16436 16804 16558
rect 17126 16532 17132 16584
rect 17184 16572 17190 16584
rect 17256 16575 17314 16581
rect 17256 16572 17268 16575
rect 17184 16544 17268 16572
rect 17184 16532 17190 16544
rect 17256 16541 17268 16544
rect 17302 16541 17314 16575
rect 17256 16535 17314 16541
rect 19978 16464 19984 16516
rect 20036 16504 20042 16516
rect 20073 16507 20131 16513
rect 20073 16504 20085 16507
rect 20036 16476 20085 16504
rect 20036 16464 20042 16476
rect 20073 16473 20085 16476
rect 20119 16504 20131 16507
rect 20162 16504 20168 16516
rect 20119 16476 20168 16504
rect 20119 16473 20131 16476
rect 20073 16467 20131 16473
rect 20162 16464 20168 16476
rect 20220 16464 20226 16516
rect 17402 16436 17408 16448
rect 16632 16408 17408 16436
rect 16632 16396 16638 16408
rect 17402 16396 17408 16408
rect 17460 16396 17466 16448
rect 1104 16346 20859 16368
rect 1104 16294 5848 16346
rect 5900 16294 5912 16346
rect 5964 16294 5976 16346
rect 6028 16294 6040 16346
rect 6092 16294 6104 16346
rect 6156 16294 10747 16346
rect 10799 16294 10811 16346
rect 10863 16294 10875 16346
rect 10927 16294 10939 16346
rect 10991 16294 11003 16346
rect 11055 16294 15646 16346
rect 15698 16294 15710 16346
rect 15762 16294 15774 16346
rect 15826 16294 15838 16346
rect 15890 16294 15902 16346
rect 15954 16294 20545 16346
rect 20597 16294 20609 16346
rect 20661 16294 20673 16346
rect 20725 16294 20737 16346
rect 20789 16294 20801 16346
rect 20853 16294 20859 16346
rect 1104 16272 20859 16294
rect 9858 16192 9864 16244
rect 9916 16192 9922 16244
rect 20070 16192 20076 16244
rect 20128 16232 20134 16244
rect 20257 16235 20315 16241
rect 20257 16232 20269 16235
rect 20128 16204 20269 16232
rect 20128 16192 20134 16204
rect 20257 16201 20269 16204
rect 20303 16201 20315 16235
rect 20257 16195 20315 16201
rect 7834 16124 7840 16176
rect 7892 16124 7898 16176
rect 17954 16124 17960 16176
rect 18012 16164 18018 16176
rect 18785 16167 18843 16173
rect 18785 16164 18797 16167
rect 18012 16136 18797 16164
rect 18012 16124 18018 16136
rect 18785 16133 18797 16136
rect 18831 16133 18843 16167
rect 18785 16127 18843 16133
rect 5905 16099 5963 16105
rect 5905 16065 5917 16099
rect 5951 16096 5963 16099
rect 6178 16096 6184 16108
rect 5951 16068 6184 16096
rect 5951 16065 5963 16068
rect 5905 16059 5963 16065
rect 6178 16056 6184 16068
rect 6236 16096 6242 16108
rect 6549 16099 6607 16105
rect 6549 16096 6561 16099
rect 6236 16068 6561 16096
rect 6236 16056 6242 16068
rect 6549 16065 6561 16068
rect 6595 16065 6607 16099
rect 6549 16059 6607 16065
rect 9677 16099 9735 16105
rect 9677 16065 9689 16099
rect 9723 16065 9735 16099
rect 9677 16059 9735 16065
rect 7101 16031 7159 16037
rect 7101 16028 7113 16031
rect 6748 16000 7113 16028
rect 6748 15969 6776 16000
rect 7101 15997 7113 16000
rect 7147 15997 7159 16031
rect 7101 15991 7159 15997
rect 7377 16031 7435 16037
rect 7377 15997 7389 16031
rect 7423 16028 7435 16031
rect 8018 16028 8024 16040
rect 7423 16000 8024 16028
rect 7423 15997 7435 16000
rect 7377 15991 7435 15997
rect 8018 15988 8024 16000
rect 8076 15988 8082 16040
rect 8849 16031 8907 16037
rect 8849 15997 8861 16031
rect 8895 16028 8907 16031
rect 9214 16028 9220 16040
rect 8895 16000 9220 16028
rect 8895 15997 8907 16000
rect 8849 15991 8907 15997
rect 9214 15988 9220 16000
rect 9272 16028 9278 16040
rect 9692 16028 9720 16059
rect 11238 16056 11244 16108
rect 11296 16096 11302 16108
rect 12161 16099 12219 16105
rect 12161 16096 12173 16099
rect 11296 16068 12173 16096
rect 11296 16056 11302 16068
rect 12161 16065 12173 16068
rect 12207 16065 12219 16099
rect 12161 16059 12219 16065
rect 19886 16056 19892 16108
rect 19944 16056 19950 16108
rect 9272 16000 9720 16028
rect 9272 15988 9278 16000
rect 18506 15988 18512 16040
rect 18564 15988 18570 16040
rect 6733 15963 6791 15969
rect 6733 15929 6745 15963
rect 6779 15929 6791 15963
rect 6733 15923 6791 15929
rect 6089 15895 6147 15901
rect 6089 15861 6101 15895
rect 6135 15892 6147 15895
rect 6362 15892 6368 15904
rect 6135 15864 6368 15892
rect 6135 15861 6147 15864
rect 6089 15855 6147 15861
rect 6362 15852 6368 15864
rect 6420 15852 6426 15904
rect 12345 15895 12403 15901
rect 12345 15861 12357 15895
rect 12391 15892 12403 15895
rect 14918 15892 14924 15904
rect 12391 15864 14924 15892
rect 12391 15861 12403 15864
rect 12345 15855 12403 15861
rect 14918 15852 14924 15864
rect 14976 15852 14982 15904
rect 1104 15802 20700 15824
rect 1104 15750 3399 15802
rect 3451 15750 3463 15802
rect 3515 15750 3527 15802
rect 3579 15750 3591 15802
rect 3643 15750 3655 15802
rect 3707 15750 8298 15802
rect 8350 15750 8362 15802
rect 8414 15750 8426 15802
rect 8478 15750 8490 15802
rect 8542 15750 8554 15802
rect 8606 15750 13197 15802
rect 13249 15750 13261 15802
rect 13313 15750 13325 15802
rect 13377 15750 13389 15802
rect 13441 15750 13453 15802
rect 13505 15750 18096 15802
rect 18148 15750 18160 15802
rect 18212 15750 18224 15802
rect 18276 15750 18288 15802
rect 18340 15750 18352 15802
rect 18404 15750 20700 15802
rect 1104 15728 20700 15750
rect 3050 15648 3056 15700
rect 3108 15688 3114 15700
rect 3191 15691 3249 15697
rect 3191 15688 3203 15691
rect 3108 15660 3203 15688
rect 3108 15648 3114 15660
rect 3191 15657 3203 15660
rect 3237 15657 3249 15691
rect 3191 15651 3249 15657
rect 3326 15648 3332 15700
rect 3384 15688 3390 15700
rect 3421 15691 3479 15697
rect 3421 15688 3433 15691
rect 3384 15660 3433 15688
rect 3384 15648 3390 15660
rect 3421 15657 3433 15660
rect 3467 15688 3479 15691
rect 3970 15688 3976 15700
rect 3467 15660 3976 15688
rect 3467 15657 3479 15660
rect 3421 15651 3479 15657
rect 3970 15648 3976 15660
rect 4028 15648 4034 15700
rect 11238 15648 11244 15700
rect 11296 15648 11302 15700
rect 13357 15691 13415 15697
rect 13357 15657 13369 15691
rect 13403 15688 13415 15691
rect 14182 15688 14188 15700
rect 13403 15660 14188 15688
rect 13403 15657 13415 15660
rect 13357 15651 13415 15657
rect 14182 15648 14188 15660
rect 14240 15648 14246 15700
rect 15378 15648 15384 15700
rect 15436 15688 15442 15700
rect 15436 15660 16620 15688
rect 15436 15648 15442 15660
rect 8573 15623 8631 15629
rect 8573 15589 8585 15623
rect 8619 15589 8631 15623
rect 14366 15620 14372 15632
rect 8573 15583 8631 15589
rect 14200 15592 14372 15620
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15552 1455 15555
rect 3234 15552 3240 15564
rect 1443 15524 3240 15552
rect 1443 15521 1455 15524
rect 1397 15515 1455 15521
rect 3234 15512 3240 15524
rect 3292 15512 3298 15564
rect 8588 15552 8616 15583
rect 8941 15555 8999 15561
rect 8941 15552 8953 15555
rect 8588 15524 8953 15552
rect 8941 15521 8953 15524
rect 8987 15521 8999 15555
rect 8941 15515 8999 15521
rect 9214 15512 9220 15564
rect 9272 15512 9278 15564
rect 11532 15524 13124 15552
rect 1762 15444 1768 15496
rect 1820 15444 1826 15496
rect 3970 15493 3976 15496
rect 3605 15487 3663 15493
rect 3605 15453 3617 15487
rect 3651 15453 3663 15487
rect 3605 15447 3663 15453
rect 3938 15487 3976 15493
rect 3938 15453 3950 15487
rect 3938 15447 3976 15453
rect 2682 15376 2688 15428
rect 2740 15376 2746 15428
rect 3620 15416 3648 15447
rect 3970 15444 3976 15447
rect 4028 15444 4034 15496
rect 4982 15444 4988 15496
rect 5040 15484 5046 15496
rect 5077 15487 5135 15493
rect 5077 15484 5089 15487
rect 5040 15456 5089 15484
rect 5040 15444 5046 15456
rect 5077 15453 5089 15456
rect 5123 15453 5135 15487
rect 5077 15447 5135 15453
rect 7009 15487 7067 15493
rect 7009 15453 7021 15487
rect 7055 15484 7067 15487
rect 7653 15487 7711 15493
rect 7653 15484 7665 15487
rect 7055 15456 7665 15484
rect 7055 15453 7067 15456
rect 7009 15447 7067 15453
rect 7653 15453 7665 15456
rect 7699 15453 7711 15487
rect 7653 15447 7711 15453
rect 7742 15444 7748 15496
rect 7800 15484 7806 15496
rect 7800 15456 8340 15484
rect 7800 15444 7806 15456
rect 7469 15419 7527 15425
rect 3620 15388 4016 15416
rect 3988 15360 4016 15388
rect 7469 15385 7481 15419
rect 7515 15416 7527 15419
rect 8312 15416 8340 15456
rect 8386 15444 8392 15496
rect 8444 15444 8450 15496
rect 11057 15487 11115 15493
rect 11057 15484 11069 15487
rect 10704 15456 11069 15484
rect 9674 15416 9680 15428
rect 7515 15388 7880 15416
rect 8312 15388 9680 15416
rect 7515 15385 7527 15388
rect 7469 15379 7527 15385
rect 3510 15308 3516 15360
rect 3568 15348 3574 15360
rect 3835 15351 3893 15357
rect 3835 15348 3847 15351
rect 3568 15320 3847 15348
rect 3568 15308 3574 15320
rect 3835 15317 3847 15320
rect 3881 15317 3893 15351
rect 3835 15311 3893 15317
rect 3970 15308 3976 15360
rect 4028 15308 4034 15360
rect 7377 15351 7435 15357
rect 7377 15317 7389 15351
rect 7423 15348 7435 15351
rect 7742 15348 7748 15360
rect 7423 15320 7748 15348
rect 7423 15317 7435 15320
rect 7377 15311 7435 15317
rect 7742 15308 7748 15320
rect 7800 15308 7806 15360
rect 7852 15357 7880 15388
rect 9674 15376 9680 15388
rect 9732 15376 9738 15428
rect 7837 15351 7895 15357
rect 7837 15317 7849 15351
rect 7883 15348 7895 15351
rect 8662 15348 8668 15360
rect 7883 15320 8668 15348
rect 7883 15317 7895 15320
rect 7837 15311 7895 15317
rect 8662 15308 8668 15320
rect 8720 15308 8726 15360
rect 9950 15308 9956 15360
rect 10008 15348 10014 15360
rect 10704 15357 10732 15456
rect 11057 15453 11069 15456
rect 11103 15453 11115 15487
rect 11057 15447 11115 15453
rect 11384 15487 11442 15493
rect 11384 15453 11396 15487
rect 11430 15484 11442 15487
rect 11532 15484 11560 15524
rect 11430 15456 11560 15484
rect 11430 15453 11442 15456
rect 11384 15447 11442 15453
rect 11606 15444 11612 15496
rect 11664 15444 11670 15496
rect 13096 15484 13124 15524
rect 14200 15493 14228 15592
rect 14366 15580 14372 15592
rect 14424 15620 14430 15632
rect 14424 15592 15056 15620
rect 14424 15580 14430 15592
rect 14918 15512 14924 15564
rect 14976 15512 14982 15564
rect 15028 15552 15056 15592
rect 15197 15555 15255 15561
rect 15197 15552 15209 15555
rect 15028 15524 15209 15552
rect 15197 15521 15209 15524
rect 15243 15552 15255 15555
rect 16592 15552 16620 15660
rect 19334 15648 19340 15700
rect 19392 15688 19398 15700
rect 19978 15688 19984 15700
rect 19392 15660 19984 15688
rect 19392 15648 19398 15660
rect 19978 15648 19984 15660
rect 20036 15688 20042 15700
rect 20073 15691 20131 15697
rect 20073 15688 20085 15691
rect 20036 15660 20085 15688
rect 20036 15648 20042 15660
rect 20073 15657 20085 15660
rect 20119 15657 20131 15691
rect 20073 15651 20131 15657
rect 16669 15623 16727 15629
rect 16669 15589 16681 15623
rect 16715 15620 16727 15623
rect 16715 15592 16896 15620
rect 16715 15589 16727 15592
rect 16669 15583 16727 15589
rect 16761 15555 16819 15561
rect 16761 15552 16773 15555
rect 15243 15524 16436 15552
rect 16592 15524 16773 15552
rect 15243 15521 15255 15524
rect 15197 15515 15255 15521
rect 13598 15487 13656 15493
rect 13598 15484 13610 15487
rect 13096 15456 13610 15484
rect 13598 15453 13610 15456
rect 13644 15484 13656 15487
rect 14160 15487 14228 15493
rect 14160 15484 14172 15487
rect 13644 15456 14172 15484
rect 13644 15453 13656 15456
rect 13598 15447 13656 15453
rect 14160 15453 14172 15456
rect 14206 15456 14228 15487
rect 16408 15484 16436 15524
rect 16761 15521 16773 15524
rect 16807 15521 16819 15555
rect 16868 15552 16896 15592
rect 17126 15552 17132 15564
rect 16868 15524 17132 15552
rect 16761 15515 16819 15521
rect 17126 15512 17132 15524
rect 17184 15512 17190 15564
rect 16408 15456 16574 15484
rect 14206 15453 14218 15456
rect 14160 15447 14218 15453
rect 11471 15419 11529 15425
rect 11471 15385 11483 15419
rect 11517 15416 11529 15419
rect 11885 15419 11943 15425
rect 11885 15416 11897 15419
rect 11517 15388 11897 15416
rect 11517 15385 11529 15388
rect 11471 15379 11529 15385
rect 11885 15385 11897 15388
rect 11931 15385 11943 15419
rect 11885 15379 11943 15385
rect 12434 15376 12440 15428
rect 12492 15376 12498 15428
rect 13262 15376 13268 15428
rect 13320 15416 13326 15428
rect 13495 15419 13553 15425
rect 13495 15416 13507 15419
rect 13320 15388 13507 15416
rect 13320 15376 13326 15388
rect 13495 15385 13507 15388
rect 13541 15385 13553 15419
rect 13495 15379 13553 15385
rect 14550 15376 14556 15428
rect 14608 15416 14614 15428
rect 16546 15416 16574 15456
rect 19794 15444 19800 15496
rect 19852 15444 19858 15496
rect 17037 15419 17095 15425
rect 17037 15416 17049 15419
rect 14608 15388 15686 15416
rect 16546 15388 17049 15416
rect 14608 15376 14614 15388
rect 14274 15357 14280 15360
rect 10689 15351 10747 15357
rect 10689 15348 10701 15351
rect 10008 15320 10701 15348
rect 10008 15308 10014 15320
rect 10689 15317 10701 15320
rect 10735 15317 10747 15351
rect 10689 15311 10747 15317
rect 14231 15351 14280 15357
rect 14231 15317 14243 15351
rect 14277 15317 14280 15351
rect 14231 15311 14280 15317
rect 14274 15308 14280 15311
rect 14332 15308 14338 15360
rect 15580 15348 15608 15388
rect 17037 15385 17049 15388
rect 17083 15385 17095 15419
rect 17494 15416 17500 15428
rect 17037 15379 17095 15385
rect 17144 15388 17500 15416
rect 17144 15348 17172 15388
rect 17494 15376 17500 15388
rect 17552 15376 17558 15428
rect 19426 15376 19432 15428
rect 19484 15416 19490 15428
rect 19981 15419 20039 15425
rect 19981 15416 19993 15419
rect 19484 15388 19993 15416
rect 19484 15376 19490 15388
rect 19981 15385 19993 15388
rect 20027 15385 20039 15419
rect 19981 15379 20039 15385
rect 15580 15320 17172 15348
rect 18506 15308 18512 15360
rect 18564 15308 18570 15360
rect 19242 15308 19248 15360
rect 19300 15348 19306 15360
rect 19613 15351 19671 15357
rect 19613 15348 19625 15351
rect 19300 15320 19625 15348
rect 19300 15308 19306 15320
rect 19613 15317 19625 15320
rect 19659 15317 19671 15351
rect 19613 15311 19671 15317
rect 1104 15258 20859 15280
rect 1104 15206 5848 15258
rect 5900 15206 5912 15258
rect 5964 15206 5976 15258
rect 6028 15206 6040 15258
rect 6092 15206 6104 15258
rect 6156 15206 10747 15258
rect 10799 15206 10811 15258
rect 10863 15206 10875 15258
rect 10927 15206 10939 15258
rect 10991 15206 11003 15258
rect 11055 15206 15646 15258
rect 15698 15206 15710 15258
rect 15762 15206 15774 15258
rect 15826 15206 15838 15258
rect 15890 15206 15902 15258
rect 15954 15206 20545 15258
rect 20597 15206 20609 15258
rect 20661 15206 20673 15258
rect 20725 15206 20737 15258
rect 20789 15206 20801 15258
rect 20853 15206 20859 15258
rect 1104 15184 20859 15206
rect 1762 15104 1768 15156
rect 1820 15144 1826 15156
rect 1903 15147 1961 15153
rect 1903 15144 1915 15147
rect 1820 15116 1915 15144
rect 1820 15104 1826 15116
rect 1903 15113 1915 15116
rect 1949 15113 1961 15147
rect 1903 15107 1961 15113
rect 2130 15104 2136 15156
rect 2188 15144 2194 15156
rect 2682 15144 2688 15156
rect 2188 15116 2688 15144
rect 2188 15104 2194 15116
rect 2682 15104 2688 15116
rect 2740 15144 2746 15156
rect 4890 15153 4896 15156
rect 4847 15147 4896 15153
rect 2740 15116 3740 15144
rect 2740 15104 2746 15116
rect 3712 15076 3740 15116
rect 4847 15113 4859 15147
rect 4893 15113 4896 15147
rect 4847 15107 4896 15113
rect 4890 15104 4896 15107
rect 4948 15104 4954 15156
rect 5997 15147 6055 15153
rect 5997 15113 6009 15147
rect 6043 15144 6055 15147
rect 6178 15144 6184 15156
rect 6043 15116 6184 15144
rect 6043 15113 6055 15116
rect 5997 15107 6055 15113
rect 6178 15104 6184 15116
rect 6236 15104 6242 15156
rect 7374 15144 7380 15156
rect 7024 15116 7380 15144
rect 7024 15076 7052 15116
rect 7374 15104 7380 15116
rect 7432 15144 7438 15156
rect 7432 15116 7972 15144
rect 7432 15104 7438 15116
rect 3712 15048 3818 15076
rect 6196 15048 7052 15076
rect 2006 15011 2064 15017
rect 2006 14977 2018 15011
rect 2052 15008 2064 15011
rect 3326 15008 3332 15020
rect 2052 14980 3332 15008
rect 2052 14977 2064 14980
rect 2006 14971 2064 14977
rect 3326 14968 3332 14980
rect 3384 14968 3390 15020
rect 3421 15011 3479 15017
rect 3421 14977 3433 15011
rect 3467 15008 3479 15011
rect 3510 15008 3516 15020
rect 3467 14980 3516 15008
rect 3467 14977 3479 14980
rect 3421 14971 3479 14977
rect 3510 14968 3516 14980
rect 3568 14968 3574 15020
rect 6196 15017 6224 15048
rect 6181 15011 6239 15017
rect 6181 14977 6193 15011
rect 6227 14977 6239 15011
rect 6181 14971 6239 14977
rect 6362 14968 6368 15020
rect 6420 14968 6426 15020
rect 7742 14968 7748 15020
rect 7800 14968 7806 15020
rect 7944 15008 7972 15116
rect 8018 15104 8024 15156
rect 8076 15144 8082 15156
rect 8113 15147 8171 15153
rect 8113 15144 8125 15147
rect 8076 15116 8125 15144
rect 8076 15104 8082 15116
rect 8113 15113 8125 15116
rect 8159 15113 8171 15147
rect 8113 15107 8171 15113
rect 8386 15104 8392 15156
rect 8444 15104 8450 15156
rect 9766 15104 9772 15156
rect 9824 15144 9830 15156
rect 11885 15147 11943 15153
rect 11885 15144 11897 15147
rect 9824 15116 10088 15144
rect 9824 15104 9830 15116
rect 8205 15011 8263 15017
rect 8205 15008 8217 15011
rect 7944 14980 8217 15008
rect 8205 14977 8217 14980
rect 8251 14977 8263 15011
rect 8404 15008 8432 15104
rect 9677 15079 9735 15085
rect 9677 15045 9689 15079
rect 9723 15076 9735 15079
rect 9950 15076 9956 15088
rect 9723 15048 9956 15076
rect 9723 15045 9735 15048
rect 9677 15039 9735 15045
rect 9950 15036 9956 15048
rect 10008 15036 10014 15088
rect 10060 15076 10088 15116
rect 11716 15116 11897 15144
rect 11716 15085 11744 15116
rect 11885 15113 11897 15116
rect 11931 15113 11943 15147
rect 11885 15107 11943 15113
rect 14737 15147 14795 15153
rect 14737 15113 14749 15147
rect 14783 15144 14795 15147
rect 15010 15144 15016 15156
rect 14783 15116 15016 15144
rect 14783 15113 14795 15116
rect 14737 15107 14795 15113
rect 15010 15104 15016 15116
rect 15068 15104 15074 15156
rect 17129 15147 17187 15153
rect 17129 15113 17141 15147
rect 17175 15144 17187 15147
rect 17954 15144 17960 15156
rect 17175 15116 17960 15144
rect 17175 15113 17187 15116
rect 17129 15107 17187 15113
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 18509 15147 18567 15153
rect 18509 15113 18521 15147
rect 18555 15113 18567 15147
rect 18509 15107 18567 15113
rect 11701 15079 11759 15085
rect 10060 15048 10166 15076
rect 11701 15045 11713 15079
rect 11747 15045 11759 15079
rect 11701 15039 11759 15045
rect 13262 15036 13268 15088
rect 13320 15036 13326 15088
rect 13998 15036 14004 15088
rect 14056 15036 14062 15088
rect 18524 15076 18552 15107
rect 19794 15104 19800 15156
rect 19852 15144 19858 15156
rect 20349 15147 20407 15153
rect 20349 15144 20361 15147
rect 19852 15116 20361 15144
rect 19852 15104 19858 15116
rect 20349 15113 20361 15116
rect 20395 15113 20407 15147
rect 20349 15107 20407 15113
rect 18877 15079 18935 15085
rect 18877 15076 18889 15079
rect 18524 15048 18889 15076
rect 18877 15045 18889 15048
rect 18923 15045 18935 15079
rect 18877 15039 18935 15045
rect 19886 15036 19892 15088
rect 19944 15036 19950 15088
rect 8665 15011 8723 15017
rect 8665 15008 8677 15011
rect 8404 14980 8677 15008
rect 8205 14971 8263 14977
rect 8665 14977 8677 14980
rect 8711 14977 8723 15011
rect 8665 14971 8723 14977
rect 11146 14968 11152 15020
rect 11204 15008 11210 15020
rect 12069 15011 12127 15017
rect 12069 15008 12081 15011
rect 11204 14980 12081 15008
rect 11204 14968 11210 14980
rect 12069 14977 12081 14980
rect 12115 14977 12127 15011
rect 18506 15008 18512 15020
rect 18354 14980 18512 15008
rect 12069 14971 12127 14977
rect 18506 14968 18512 14980
rect 18564 14968 18570 15020
rect 3050 14900 3056 14952
rect 3108 14900 3114 14952
rect 5166 14900 5172 14952
rect 5224 14940 5230 14952
rect 6641 14943 6699 14949
rect 6641 14940 6653 14943
rect 5224 14912 6653 14940
rect 5224 14900 5230 14912
rect 6641 14909 6653 14912
rect 6687 14909 6699 14943
rect 6641 14903 6699 14909
rect 9401 14943 9459 14949
rect 9401 14909 9413 14943
rect 9447 14909 9459 14943
rect 9401 14903 9459 14909
rect 11517 14943 11575 14949
rect 11517 14909 11529 14943
rect 11563 14940 11575 14943
rect 11606 14940 11612 14952
rect 11563 14912 11612 14940
rect 11563 14909 11575 14912
rect 11517 14903 11575 14909
rect 8849 14875 8907 14881
rect 8849 14841 8861 14875
rect 8895 14872 8907 14875
rect 9416 14872 9444 14903
rect 11606 14900 11612 14912
rect 11664 14940 11670 14952
rect 12989 14943 13047 14949
rect 12989 14940 13001 14943
rect 11664 14912 13001 14940
rect 11664 14900 11670 14912
rect 12989 14909 13001 14912
rect 13035 14940 13047 14943
rect 13906 14940 13912 14952
rect 13035 14912 13912 14940
rect 13035 14909 13047 14912
rect 12989 14903 13047 14909
rect 13906 14900 13912 14912
rect 13964 14900 13970 14952
rect 17678 14900 17684 14952
rect 17736 14900 17742 14952
rect 18598 14900 18604 14952
rect 18656 14900 18662 14952
rect 8895 14844 9444 14872
rect 8895 14841 8907 14844
rect 8849 14835 8907 14841
rect 17034 14832 17040 14884
rect 17092 14872 17098 14884
rect 18141 14875 18199 14881
rect 18141 14872 18153 14875
rect 17092 14844 18153 14872
rect 17092 14832 17098 14844
rect 18141 14841 18153 14844
rect 18187 14841 18199 14875
rect 18141 14835 18199 14841
rect 11146 14764 11152 14816
rect 11204 14764 11210 14816
rect 1104 14714 20700 14736
rect 1104 14662 3399 14714
rect 3451 14662 3463 14714
rect 3515 14662 3527 14714
rect 3579 14662 3591 14714
rect 3643 14662 3655 14714
rect 3707 14662 8298 14714
rect 8350 14662 8362 14714
rect 8414 14662 8426 14714
rect 8478 14662 8490 14714
rect 8542 14662 8554 14714
rect 8606 14662 13197 14714
rect 13249 14662 13261 14714
rect 13313 14662 13325 14714
rect 13377 14662 13389 14714
rect 13441 14662 13453 14714
rect 13505 14662 18096 14714
rect 18148 14662 18160 14714
rect 18212 14662 18224 14714
rect 18276 14662 18288 14714
rect 18340 14662 18352 14714
rect 18404 14662 20700 14714
rect 1104 14640 20700 14662
rect 5166 14560 5172 14612
rect 5224 14560 5230 14612
rect 15841 14603 15899 14609
rect 15841 14569 15853 14603
rect 15887 14600 15899 14603
rect 16574 14600 16580 14612
rect 15887 14572 16580 14600
rect 15887 14569 15899 14572
rect 15841 14563 15899 14569
rect 16574 14560 16580 14572
rect 16632 14560 16638 14612
rect 17034 14560 17040 14612
rect 17092 14560 17098 14612
rect 17218 14492 17224 14544
rect 17276 14532 17282 14544
rect 18049 14535 18107 14541
rect 18049 14532 18061 14535
rect 17276 14504 18061 14532
rect 17276 14492 17282 14504
rect 18049 14501 18061 14504
rect 18095 14501 18107 14535
rect 18049 14495 18107 14501
rect 13906 14424 13912 14476
rect 13964 14464 13970 14476
rect 14093 14467 14151 14473
rect 14093 14464 14105 14467
rect 13964 14436 14105 14464
rect 13964 14424 13970 14436
rect 14093 14433 14105 14436
rect 14139 14433 14151 14467
rect 14093 14427 14151 14433
rect 17678 14424 17684 14476
rect 17736 14424 17742 14476
rect 4982 14356 4988 14408
rect 5040 14356 5046 14408
rect 17126 14356 17132 14408
rect 17184 14396 17190 14408
rect 17184 14368 17250 14396
rect 17184 14356 17190 14368
rect 14274 14288 14280 14340
rect 14332 14328 14338 14340
rect 14369 14331 14427 14337
rect 14369 14328 14381 14331
rect 14332 14300 14381 14328
rect 14332 14288 14338 14300
rect 14369 14297 14381 14300
rect 14415 14297 14427 14331
rect 14369 14291 14427 14297
rect 15378 14288 15384 14340
rect 15436 14288 15442 14340
rect 18414 14220 18420 14272
rect 18472 14220 18478 14272
rect 1104 14170 20859 14192
rect 1104 14118 5848 14170
rect 5900 14118 5912 14170
rect 5964 14118 5976 14170
rect 6028 14118 6040 14170
rect 6092 14118 6104 14170
rect 6156 14118 10747 14170
rect 10799 14118 10811 14170
rect 10863 14118 10875 14170
rect 10927 14118 10939 14170
rect 10991 14118 11003 14170
rect 11055 14118 15646 14170
rect 15698 14118 15710 14170
rect 15762 14118 15774 14170
rect 15826 14118 15838 14170
rect 15890 14118 15902 14170
rect 15954 14118 20545 14170
rect 20597 14118 20609 14170
rect 20661 14118 20673 14170
rect 20725 14118 20737 14170
rect 20789 14118 20801 14170
rect 20853 14118 20859 14170
rect 1104 14096 20859 14118
rect 8662 13948 8668 14000
rect 8720 13948 8726 14000
rect 18414 13948 18420 14000
rect 18472 13988 18478 14000
rect 18877 13991 18935 13997
rect 18877 13988 18889 13991
rect 18472 13960 18889 13988
rect 18472 13948 18478 13960
rect 18877 13957 18889 13960
rect 18923 13957 18935 13991
rect 18877 13951 18935 13957
rect 19886 13948 19892 14000
rect 19944 13948 19950 14000
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 2222 13880 2228 13932
rect 2280 13880 2286 13932
rect 13078 13880 13084 13932
rect 13136 13920 13142 13932
rect 13300 13923 13358 13929
rect 13300 13920 13312 13923
rect 13136 13892 13312 13920
rect 13136 13880 13142 13892
rect 13300 13889 13312 13892
rect 13346 13889 13358 13923
rect 13300 13883 13358 13889
rect 14093 13923 14151 13929
rect 14093 13889 14105 13923
rect 14139 13920 14151 13923
rect 14550 13920 14556 13932
rect 14139 13892 14556 13920
rect 14139 13889 14151 13892
rect 14093 13883 14151 13889
rect 3970 13812 3976 13864
rect 4028 13812 4034 13864
rect 7834 13812 7840 13864
rect 7892 13812 7898 13864
rect 13403 13855 13461 13861
rect 13403 13821 13415 13855
rect 13449 13852 13461 13855
rect 13909 13855 13967 13861
rect 13909 13852 13921 13855
rect 13449 13824 13921 13852
rect 13449 13821 13461 13824
rect 13403 13815 13461 13821
rect 13909 13821 13921 13824
rect 13955 13821 13967 13855
rect 13909 13815 13967 13821
rect 11146 13784 11152 13796
rect 9508 13756 11152 13784
rect 1486 13676 1492 13728
rect 1544 13716 1550 13728
rect 1581 13719 1639 13725
rect 1581 13716 1593 13719
rect 1544 13688 1593 13716
rect 1544 13676 1550 13688
rect 1581 13685 1593 13688
rect 1627 13685 1639 13719
rect 1581 13679 1639 13685
rect 8100 13719 8158 13725
rect 8100 13685 8112 13719
rect 8146 13716 8158 13719
rect 9508 13716 9536 13756
rect 11146 13744 11152 13756
rect 11204 13744 11210 13796
rect 12526 13744 12532 13796
rect 12584 13784 12590 13796
rect 14108 13784 14136 13883
rect 14550 13880 14556 13892
rect 14608 13880 14614 13932
rect 14277 13855 14335 13861
rect 14277 13821 14289 13855
rect 14323 13852 14335 13855
rect 15378 13852 15384 13864
rect 14323 13824 15384 13852
rect 14323 13821 14335 13824
rect 14277 13815 14335 13821
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 18598 13812 18604 13864
rect 18656 13812 18662 13864
rect 12584 13756 14136 13784
rect 12584 13744 12590 13756
rect 8146 13688 9536 13716
rect 8146 13685 8158 13688
rect 8100 13679 8158 13685
rect 9582 13676 9588 13728
rect 9640 13676 9646 13728
rect 20346 13676 20352 13728
rect 20404 13676 20410 13728
rect 1104 13626 20700 13648
rect 1104 13574 3399 13626
rect 3451 13574 3463 13626
rect 3515 13574 3527 13626
rect 3579 13574 3591 13626
rect 3643 13574 3655 13626
rect 3707 13574 8298 13626
rect 8350 13574 8362 13626
rect 8414 13574 8426 13626
rect 8478 13574 8490 13626
rect 8542 13574 8554 13626
rect 8606 13574 13197 13626
rect 13249 13574 13261 13626
rect 13313 13574 13325 13626
rect 13377 13574 13389 13626
rect 13441 13574 13453 13626
rect 13505 13574 18096 13626
rect 18148 13574 18160 13626
rect 18212 13574 18224 13626
rect 18276 13574 18288 13626
rect 18340 13574 18352 13626
rect 18404 13574 20700 13626
rect 1104 13552 20700 13574
rect 7834 13472 7840 13524
rect 7892 13472 7898 13524
rect 10502 13472 10508 13524
rect 10560 13512 10566 13524
rect 12253 13515 12311 13521
rect 12253 13512 12265 13515
rect 10560 13484 12265 13512
rect 10560 13472 10566 13484
rect 12253 13481 12265 13484
rect 12299 13481 12311 13515
rect 12253 13475 12311 13481
rect 13078 13472 13084 13524
rect 13136 13472 13142 13524
rect 17402 13472 17408 13524
rect 17460 13472 17466 13524
rect 1673 13447 1731 13453
rect 1673 13413 1685 13447
rect 1719 13413 1731 13447
rect 1673 13407 1731 13413
rect 7561 13447 7619 13453
rect 7561 13413 7573 13447
rect 7607 13413 7619 13447
rect 7561 13407 7619 13413
rect 9953 13447 10011 13453
rect 9953 13413 9965 13447
rect 9999 13444 10011 13447
rect 12526 13444 12532 13456
rect 9999 13416 10456 13444
rect 9999 13413 10011 13416
rect 9953 13407 10011 13413
rect 1486 13268 1492 13320
rect 1544 13268 1550 13320
rect 1688 13308 1716 13407
rect 2222 13336 2228 13388
rect 2280 13336 2286 13388
rect 1857 13311 1915 13317
rect 1857 13308 1869 13311
rect 1688 13280 1869 13308
rect 1857 13277 1869 13280
rect 1903 13277 1915 13311
rect 1857 13271 1915 13277
rect 4890 13268 4896 13320
rect 4948 13308 4954 13320
rect 4985 13311 5043 13317
rect 4985 13308 4997 13311
rect 4948 13280 4997 13308
rect 4948 13268 4954 13280
rect 4985 13277 4997 13280
rect 5031 13277 5043 13311
rect 5445 13311 5503 13317
rect 5445 13308 5457 13311
rect 4985 13271 5043 13277
rect 5184 13280 5457 13308
rect 5184 13181 5212 13280
rect 5445 13277 5457 13280
rect 5491 13277 5503 13311
rect 5445 13271 5503 13277
rect 7374 13268 7380 13320
rect 7432 13268 7438 13320
rect 7576 13308 7604 13407
rect 10428 13320 10456 13416
rect 11808 13416 12532 13444
rect 7653 13311 7711 13317
rect 7653 13308 7665 13311
rect 7576 13280 7665 13308
rect 7653 13277 7665 13280
rect 7699 13308 7711 13311
rect 7834 13308 7840 13320
rect 7699 13280 7840 13308
rect 7699 13277 7711 13280
rect 7653 13271 7711 13277
rect 7834 13268 7840 13280
rect 7892 13268 7898 13320
rect 8478 13268 8484 13320
rect 8536 13308 8542 13320
rect 9493 13311 9551 13317
rect 9493 13308 9505 13311
rect 8536 13280 9505 13308
rect 8536 13268 8542 13280
rect 9493 13277 9505 13280
rect 9539 13308 9551 13311
rect 9582 13308 9588 13320
rect 9539 13280 9588 13308
rect 9539 13277 9551 13280
rect 9493 13271 9551 13277
rect 9582 13268 9588 13280
rect 9640 13268 9646 13320
rect 9769 13311 9827 13317
rect 9769 13308 9781 13311
rect 9692 13280 9781 13308
rect 5169 13175 5227 13181
rect 5169 13141 5181 13175
rect 5215 13141 5227 13175
rect 5169 13135 5227 13141
rect 5629 13175 5687 13181
rect 5629 13141 5641 13175
rect 5675 13172 5687 13175
rect 6914 13172 6920 13184
rect 5675 13144 6920 13172
rect 5675 13141 5687 13144
rect 5629 13135 5687 13141
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 9692 13181 9720 13280
rect 9769 13277 9781 13280
rect 9815 13277 9827 13311
rect 9769 13271 9827 13277
rect 9858 13268 9864 13320
rect 9916 13308 9922 13320
rect 10045 13311 10103 13317
rect 10045 13308 10057 13311
rect 9916 13280 10057 13308
rect 9916 13268 9922 13280
rect 10045 13277 10057 13280
rect 10091 13277 10103 13311
rect 10045 13271 10103 13277
rect 10410 13268 10416 13320
rect 10468 13268 10474 13320
rect 11808 13294 11836 13416
rect 12526 13404 12532 13416
rect 12584 13404 12590 13456
rect 20162 13404 20168 13456
rect 20220 13404 20226 13456
rect 12158 13336 12164 13388
rect 12216 13376 12222 13388
rect 12713 13379 12771 13385
rect 12713 13376 12725 13379
rect 12216 13348 12725 13376
rect 12216 13336 12222 13348
rect 12713 13345 12725 13348
rect 12759 13345 12771 13379
rect 12713 13339 12771 13345
rect 13906 13336 13912 13388
rect 13964 13376 13970 13388
rect 14093 13379 14151 13385
rect 14093 13376 14105 13379
rect 13964 13348 14105 13376
rect 13964 13336 13970 13348
rect 14093 13345 14105 13348
rect 14139 13345 14151 13379
rect 14093 13339 14151 13345
rect 14366 13336 14372 13388
rect 14424 13336 14430 13388
rect 11974 13268 11980 13320
rect 12032 13308 12038 13320
rect 12437 13311 12495 13317
rect 12437 13308 12449 13311
rect 12032 13280 12449 13308
rect 12032 13268 12038 13280
rect 12437 13277 12449 13280
rect 12483 13277 12495 13311
rect 12437 13271 12495 13277
rect 10594 13200 10600 13252
rect 10652 13240 10658 13252
rect 10689 13243 10747 13249
rect 10689 13240 10701 13243
rect 10652 13212 10701 13240
rect 10652 13200 10658 13212
rect 10689 13209 10701 13212
rect 10735 13209 10747 13243
rect 12452 13240 12480 13271
rect 12526 13268 12532 13320
rect 12584 13268 12590 13320
rect 12897 13311 12955 13317
rect 12897 13277 12909 13311
rect 12943 13277 12955 13311
rect 12897 13271 12955 13277
rect 12912 13240 12940 13271
rect 17402 13268 17408 13320
rect 17460 13308 17466 13320
rect 17865 13311 17923 13317
rect 17865 13308 17877 13311
rect 17460 13280 17877 13308
rect 17460 13268 17466 13280
rect 17865 13277 17877 13280
rect 17911 13277 17923 13311
rect 17865 13271 17923 13277
rect 20346 13268 20352 13320
rect 20404 13268 20410 13320
rect 12452 13212 12940 13240
rect 10689 13203 10747 13209
rect 15378 13200 15384 13252
rect 15436 13200 15442 13252
rect 16574 13200 16580 13252
rect 16632 13240 16638 13252
rect 17313 13243 17371 13249
rect 17313 13240 17325 13243
rect 16632 13212 17325 13240
rect 16632 13200 16638 13212
rect 17313 13209 17325 13212
rect 17359 13240 17371 13243
rect 18966 13240 18972 13252
rect 17359 13212 18972 13240
rect 17359 13209 17371 13212
rect 17313 13203 17371 13209
rect 18966 13200 18972 13212
rect 19024 13200 19030 13252
rect 9677 13175 9735 13181
rect 9677 13141 9689 13175
rect 9723 13141 9735 13175
rect 9677 13135 9735 13141
rect 10229 13175 10287 13181
rect 10229 13141 10241 13175
rect 10275 13172 10287 13175
rect 10318 13172 10324 13184
rect 10275 13144 10324 13172
rect 10275 13141 10287 13144
rect 10229 13135 10287 13141
rect 10318 13132 10324 13144
rect 10376 13132 10382 13184
rect 15841 13175 15899 13181
rect 15841 13141 15853 13175
rect 15887 13172 15899 13175
rect 16022 13172 16028 13184
rect 15887 13144 16028 13172
rect 15887 13141 15899 13144
rect 15841 13135 15899 13141
rect 16022 13132 16028 13144
rect 16080 13132 16086 13184
rect 18046 13132 18052 13184
rect 18104 13172 18110 13184
rect 18141 13175 18199 13181
rect 18141 13172 18153 13175
rect 18104 13144 18153 13172
rect 18104 13132 18110 13144
rect 18141 13141 18153 13144
rect 18187 13141 18199 13175
rect 18141 13135 18199 13141
rect 1104 13082 20859 13104
rect 1104 13030 5848 13082
rect 5900 13030 5912 13082
rect 5964 13030 5976 13082
rect 6028 13030 6040 13082
rect 6092 13030 6104 13082
rect 6156 13030 10747 13082
rect 10799 13030 10811 13082
rect 10863 13030 10875 13082
rect 10927 13030 10939 13082
rect 10991 13030 11003 13082
rect 11055 13030 15646 13082
rect 15698 13030 15710 13082
rect 15762 13030 15774 13082
rect 15826 13030 15838 13082
rect 15890 13030 15902 13082
rect 15954 13030 20545 13082
rect 20597 13030 20609 13082
rect 20661 13030 20673 13082
rect 20725 13030 20737 13082
rect 20789 13030 20801 13082
rect 20853 13030 20859 13082
rect 1104 13008 20859 13030
rect 4890 12928 4896 12980
rect 4948 12928 4954 12980
rect 4985 12971 5043 12977
rect 4985 12937 4997 12971
rect 5031 12937 5043 12971
rect 4985 12931 5043 12937
rect 7009 12971 7067 12977
rect 7009 12937 7021 12971
rect 7055 12968 7067 12971
rect 7374 12968 7380 12980
rect 7055 12940 7380 12968
rect 7055 12937 7067 12940
rect 7009 12931 7067 12937
rect 4709 12835 4767 12841
rect 4709 12801 4721 12835
rect 4755 12832 4767 12835
rect 5000 12832 5028 12931
rect 7374 12928 7380 12940
rect 7432 12928 7438 12980
rect 8662 12928 8668 12980
rect 8720 12928 8726 12980
rect 11333 12971 11391 12977
rect 11333 12937 11345 12971
rect 11379 12937 11391 12971
rect 11333 12931 11391 12937
rect 8478 12860 8484 12912
rect 8536 12860 8542 12912
rect 8680 12900 8708 12928
rect 8938 12900 8944 12912
rect 8680 12872 8944 12900
rect 8938 12860 8944 12872
rect 8996 12860 9002 12912
rect 4755 12804 5028 12832
rect 4755 12801 4767 12804
rect 4709 12795 4767 12801
rect 5166 12792 5172 12844
rect 5224 12792 5230 12844
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12832 6883 12835
rect 6914 12832 6920 12844
rect 6871 12804 6920 12832
rect 6871 12801 6883 12804
rect 6825 12795 6883 12801
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 7834 12792 7840 12844
rect 7892 12792 7898 12844
rect 10226 12792 10232 12844
rect 10284 12792 10290 12844
rect 10410 12792 10416 12844
rect 10468 12832 10474 12844
rect 11149 12835 11207 12841
rect 11149 12832 11161 12835
rect 10468 12804 11161 12832
rect 10468 12792 10474 12804
rect 11149 12801 11161 12804
rect 11195 12801 11207 12835
rect 11348 12832 11376 12931
rect 11974 12928 11980 12980
rect 12032 12928 12038 12980
rect 12207 12971 12265 12977
rect 12207 12937 12219 12971
rect 12253 12968 12265 12971
rect 12526 12968 12532 12980
rect 12253 12940 12532 12968
rect 12253 12937 12265 12940
rect 12207 12931 12265 12937
rect 12526 12928 12532 12940
rect 12584 12928 12590 12980
rect 14550 12928 14556 12980
rect 14608 12968 14614 12980
rect 15102 12968 15108 12980
rect 14608 12940 15108 12968
rect 14608 12928 14614 12940
rect 15102 12928 15108 12940
rect 15160 12968 15166 12980
rect 15160 12940 18092 12968
rect 15160 12928 15166 12940
rect 12406 12872 16574 12900
rect 12158 12841 12164 12844
rect 11793 12835 11851 12841
rect 11793 12832 11805 12835
rect 11348 12804 11805 12832
rect 11149 12795 11207 12801
rect 11793 12801 11805 12804
rect 11839 12801 11851 12835
rect 11793 12795 11851 12801
rect 12136 12835 12164 12841
rect 12136 12801 12148 12835
rect 12136 12795 12164 12801
rect 8205 12767 8263 12773
rect 8205 12733 8217 12767
rect 8251 12733 8263 12767
rect 8205 12727 8263 12733
rect 8021 12699 8079 12705
rect 8021 12665 8033 12699
rect 8067 12696 8079 12699
rect 8220 12696 8248 12727
rect 10318 12724 10324 12776
rect 10376 12724 10382 12776
rect 10594 12724 10600 12776
rect 10652 12724 10658 12776
rect 11164 12764 11192 12795
rect 12158 12792 12164 12795
rect 12216 12792 12222 12844
rect 12406 12764 12434 12872
rect 16546 12832 16574 12872
rect 18064 12844 18092 12940
rect 16669 12835 16727 12841
rect 16669 12832 16681 12835
rect 16546 12804 16681 12832
rect 16669 12801 16681 12804
rect 16715 12801 16727 12835
rect 16669 12795 16727 12801
rect 18046 12792 18052 12844
rect 18104 12792 18110 12844
rect 16945 12767 17003 12773
rect 16945 12764 16957 12767
rect 11164 12736 12434 12764
rect 16776 12736 16957 12764
rect 8067 12668 8248 12696
rect 10336 12696 10364 12724
rect 11054 12696 11060 12708
rect 10336 12668 11060 12696
rect 8067 12665 8079 12668
rect 8021 12659 8079 12665
rect 11054 12656 11060 12668
rect 11112 12656 11118 12708
rect 14366 12656 14372 12708
rect 14424 12696 14430 12708
rect 14642 12696 14648 12708
rect 14424 12668 14648 12696
rect 14424 12656 14430 12668
rect 14642 12656 14648 12668
rect 14700 12696 14706 12708
rect 16776 12696 16804 12736
rect 16945 12733 16957 12736
rect 16991 12733 17003 12767
rect 16945 12727 17003 12733
rect 14700 12668 16804 12696
rect 14700 12656 14706 12668
rect 9858 12588 9864 12640
rect 9916 12628 9922 12640
rect 9953 12631 10011 12637
rect 9953 12628 9965 12631
rect 9916 12600 9965 12628
rect 9916 12588 9922 12600
rect 9953 12597 9965 12600
rect 9999 12597 10011 12631
rect 9953 12591 10011 12597
rect 18414 12588 18420 12640
rect 18472 12588 18478 12640
rect 1104 12538 20700 12560
rect 1104 12486 3399 12538
rect 3451 12486 3463 12538
rect 3515 12486 3527 12538
rect 3579 12486 3591 12538
rect 3643 12486 3655 12538
rect 3707 12486 8298 12538
rect 8350 12486 8362 12538
rect 8414 12486 8426 12538
rect 8478 12486 8490 12538
rect 8542 12486 8554 12538
rect 8606 12486 13197 12538
rect 13249 12486 13261 12538
rect 13313 12486 13325 12538
rect 13377 12486 13389 12538
rect 13441 12486 13453 12538
rect 13505 12486 18096 12538
rect 18148 12486 18160 12538
rect 18212 12486 18224 12538
rect 18276 12486 18288 12538
rect 18340 12486 18352 12538
rect 18404 12486 20700 12538
rect 1104 12464 20700 12486
rect 4709 12427 4767 12433
rect 4709 12393 4721 12427
rect 4755 12424 4767 12427
rect 5166 12424 5172 12436
rect 4755 12396 5172 12424
rect 4755 12393 4767 12396
rect 4709 12387 4767 12393
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 11054 12384 11060 12436
rect 11112 12424 11118 12436
rect 11958 12427 12016 12433
rect 11958 12424 11970 12427
rect 11112 12396 11970 12424
rect 11112 12384 11118 12396
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12220 4583 12223
rect 4571 12192 4844 12220
rect 4571 12189 4583 12192
rect 4525 12183 4583 12189
rect 4816 12093 4844 12192
rect 4982 12180 4988 12232
rect 5040 12180 5046 12232
rect 6365 12223 6423 12229
rect 6365 12189 6377 12223
rect 6411 12220 6423 12223
rect 7374 12220 7380 12232
rect 6411 12192 7380 12220
rect 6411 12189 6423 12192
rect 6365 12183 6423 12189
rect 7374 12180 7380 12192
rect 7432 12180 7438 12232
rect 4801 12087 4859 12093
rect 4801 12053 4813 12087
rect 4847 12053 4859 12087
rect 4801 12047 4859 12053
rect 6178 12044 6184 12096
rect 6236 12044 6242 12096
rect 11624 12084 11652 12396
rect 11958 12393 11970 12396
rect 12004 12393 12016 12427
rect 11958 12387 12016 12393
rect 17218 12384 17224 12436
rect 17276 12384 17282 12436
rect 16390 12316 16396 12368
rect 16448 12356 16454 12368
rect 16448 12328 17540 12356
rect 16448 12316 16454 12328
rect 11701 12291 11759 12297
rect 11701 12257 11713 12291
rect 11747 12288 11759 12291
rect 13906 12288 13912 12300
rect 11747 12260 13912 12288
rect 11747 12257 11759 12260
rect 11701 12251 11759 12257
rect 13906 12248 13912 12260
rect 13964 12288 13970 12300
rect 14369 12291 14427 12297
rect 14369 12288 14381 12291
rect 13964 12260 14381 12288
rect 13964 12248 13970 12260
rect 14369 12257 14381 12260
rect 14415 12257 14427 12291
rect 14369 12251 14427 12257
rect 14642 12248 14648 12300
rect 14700 12248 14706 12300
rect 17512 12274 17540 12328
rect 17586 12316 17592 12368
rect 17644 12356 17650 12368
rect 18233 12359 18291 12365
rect 18233 12356 18245 12359
rect 17644 12328 18245 12356
rect 17644 12316 17650 12328
rect 18233 12325 18245 12328
rect 18279 12325 18291 12359
rect 18233 12319 18291 12325
rect 18414 12180 18420 12232
rect 18472 12180 18478 12232
rect 20346 12180 20352 12232
rect 20404 12180 20410 12232
rect 12434 12112 12440 12164
rect 12492 12112 12498 12164
rect 14642 12152 14648 12164
rect 13280 12124 14648 12152
rect 13280 12084 13308 12124
rect 14642 12112 14648 12124
rect 14700 12112 14706 12164
rect 15102 12112 15108 12164
rect 15160 12112 15166 12164
rect 16390 12112 16396 12164
rect 16448 12112 16454 12164
rect 11624 12056 13308 12084
rect 13449 12087 13507 12093
rect 13449 12053 13461 12087
rect 13495 12084 13507 12087
rect 13630 12084 13636 12096
rect 13495 12056 13636 12084
rect 13495 12053 13507 12056
rect 13449 12047 13507 12053
rect 13630 12044 13636 12056
rect 13688 12044 13694 12096
rect 18601 12087 18659 12093
rect 18601 12053 18613 12087
rect 18647 12084 18659 12087
rect 18874 12084 18880 12096
rect 18647 12056 18880 12084
rect 18647 12053 18659 12056
rect 18601 12047 18659 12053
rect 18874 12044 18880 12056
rect 18932 12044 18938 12096
rect 20162 12044 20168 12096
rect 20220 12044 20226 12096
rect 1104 11994 20859 12016
rect 1104 11942 5848 11994
rect 5900 11942 5912 11994
rect 5964 11942 5976 11994
rect 6028 11942 6040 11994
rect 6092 11942 6104 11994
rect 6156 11942 10747 11994
rect 10799 11942 10811 11994
rect 10863 11942 10875 11994
rect 10927 11942 10939 11994
rect 10991 11942 11003 11994
rect 11055 11942 15646 11994
rect 15698 11942 15710 11994
rect 15762 11942 15774 11994
rect 15826 11942 15838 11994
rect 15890 11942 15902 11994
rect 15954 11942 20545 11994
rect 20597 11942 20609 11994
rect 20661 11942 20673 11994
rect 20725 11942 20737 11994
rect 20789 11942 20801 11994
rect 20853 11942 20859 11994
rect 1104 11920 20859 11942
rect 2593 11883 2651 11889
rect 2593 11849 2605 11883
rect 2639 11849 2651 11883
rect 2593 11843 2651 11849
rect 3697 11883 3755 11889
rect 3697 11849 3709 11883
rect 3743 11849 3755 11883
rect 3697 11843 3755 11849
rect 4157 11883 4215 11889
rect 4157 11849 4169 11883
rect 4203 11880 4215 11883
rect 4982 11880 4988 11892
rect 4203 11852 4988 11880
rect 4203 11849 4215 11852
rect 4157 11843 4215 11849
rect 2608 11812 2636 11843
rect 2608 11784 3004 11812
rect 1486 11704 1492 11756
rect 1544 11744 1550 11756
rect 2976 11753 3004 11784
rect 1857 11747 1915 11753
rect 1857 11744 1869 11747
rect 1544 11716 1869 11744
rect 1544 11704 1550 11716
rect 1857 11713 1869 11716
rect 1903 11713 1915 11747
rect 1857 11707 1915 11713
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11744 2467 11747
rect 2869 11747 2927 11753
rect 2455 11716 2728 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 1762 11636 1768 11688
rect 1820 11636 1826 11688
rect 2700 11617 2728 11716
rect 2869 11713 2881 11747
rect 2915 11713 2927 11747
rect 2869 11707 2927 11713
rect 2961 11747 3019 11753
rect 2961 11713 2973 11747
rect 3007 11713 3019 11747
rect 3513 11747 3571 11753
rect 3513 11744 3525 11747
rect 2961 11707 3019 11713
rect 3160 11716 3525 11744
rect 2685 11611 2743 11617
rect 2685 11577 2697 11611
rect 2731 11577 2743 11611
rect 2685 11571 2743 11577
rect 2225 11543 2283 11549
rect 2225 11509 2237 11543
rect 2271 11540 2283 11543
rect 2884 11540 2912 11707
rect 3160 11617 3188 11716
rect 3513 11713 3525 11716
rect 3559 11713 3571 11747
rect 3712 11744 3740 11843
rect 4982 11840 4988 11852
rect 5040 11840 5046 11892
rect 12069 11883 12127 11889
rect 12069 11849 12081 11883
rect 12115 11880 12127 11883
rect 12434 11880 12440 11892
rect 12115 11852 12440 11880
rect 12115 11849 12127 11852
rect 12069 11843 12127 11849
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 13814 11840 13820 11892
rect 13872 11840 13878 11892
rect 20346 11840 20352 11892
rect 20404 11840 20410 11892
rect 13832 11812 13860 11840
rect 13188 11784 13860 11812
rect 3973 11747 4031 11753
rect 3973 11744 3985 11747
rect 3712 11716 3985 11744
rect 3513 11707 3571 11713
rect 3973 11713 3985 11716
rect 4019 11713 4031 11747
rect 3973 11707 4031 11713
rect 5997 11747 6055 11753
rect 5997 11713 6009 11747
rect 6043 11744 6055 11747
rect 6178 11744 6184 11756
rect 6043 11716 6184 11744
rect 6043 11713 6055 11716
rect 5997 11707 6055 11713
rect 6178 11704 6184 11716
rect 6236 11704 6242 11756
rect 11882 11704 11888 11756
rect 11940 11704 11946 11756
rect 13188 11753 13216 11784
rect 13998 11772 14004 11824
rect 14056 11772 14062 11824
rect 18874 11772 18880 11824
rect 18932 11772 18938 11824
rect 19426 11772 19432 11824
rect 19484 11772 19490 11824
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 11698 11636 11704 11688
rect 11756 11636 11762 11688
rect 11790 11636 11796 11688
rect 11848 11676 11854 11688
rect 13449 11679 13507 11685
rect 13449 11676 13461 11679
rect 11848 11648 13461 11676
rect 11848 11636 11854 11648
rect 13449 11645 13461 11648
rect 13495 11676 13507 11679
rect 15654 11676 15660 11688
rect 13495 11648 15660 11676
rect 13495 11645 13507 11648
rect 13449 11639 13507 11645
rect 15654 11636 15660 11648
rect 15712 11636 15718 11688
rect 16206 11636 16212 11688
rect 16264 11676 16270 11688
rect 18601 11679 18659 11685
rect 18601 11676 18613 11679
rect 16264 11648 18613 11676
rect 16264 11636 16270 11648
rect 18601 11645 18613 11648
rect 18647 11645 18659 11679
rect 18601 11639 18659 11645
rect 3145 11611 3203 11617
rect 3145 11577 3157 11611
rect 3191 11577 3203 11611
rect 3145 11571 3203 11577
rect 2271 11512 2912 11540
rect 2271 11509 2283 11512
rect 2225 11503 2283 11509
rect 6178 11500 6184 11552
rect 6236 11500 6242 11552
rect 14921 11543 14979 11549
rect 14921 11509 14933 11543
rect 14967 11540 14979 11543
rect 15010 11540 15016 11552
rect 14967 11512 15016 11540
rect 14967 11509 14979 11512
rect 14921 11503 14979 11509
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 1104 11450 20700 11472
rect 1104 11398 3399 11450
rect 3451 11398 3463 11450
rect 3515 11398 3527 11450
rect 3579 11398 3591 11450
rect 3643 11398 3655 11450
rect 3707 11398 8298 11450
rect 8350 11398 8362 11450
rect 8414 11398 8426 11450
rect 8478 11398 8490 11450
rect 8542 11398 8554 11450
rect 8606 11398 13197 11450
rect 13249 11398 13261 11450
rect 13313 11398 13325 11450
rect 13377 11398 13389 11450
rect 13441 11398 13453 11450
rect 13505 11398 18096 11450
rect 18148 11398 18160 11450
rect 18212 11398 18224 11450
rect 18276 11398 18288 11450
rect 18340 11398 18352 11450
rect 18404 11398 20700 11450
rect 1104 11376 20700 11398
rect 8938 11296 8944 11348
rect 8996 11336 9002 11348
rect 9490 11336 9496 11348
rect 8996 11308 9496 11336
rect 8996 11296 9002 11308
rect 9490 11296 9496 11308
rect 9548 11336 9554 11348
rect 9585 11339 9643 11345
rect 9585 11336 9597 11339
rect 9548 11308 9597 11336
rect 9548 11296 9554 11308
rect 9585 11305 9597 11308
rect 9631 11305 9643 11339
rect 9585 11299 9643 11305
rect 11195 11339 11253 11345
rect 11195 11305 11207 11339
rect 11241 11336 11253 11339
rect 11698 11336 11704 11348
rect 11241 11308 11704 11336
rect 11241 11305 11253 11308
rect 11195 11299 11253 11305
rect 11698 11296 11704 11308
rect 11756 11296 11762 11348
rect 13998 11296 14004 11348
rect 14056 11336 14062 11348
rect 14461 11339 14519 11345
rect 14461 11336 14473 11339
rect 14056 11308 14473 11336
rect 14056 11296 14062 11308
rect 14461 11305 14473 11308
rect 14507 11305 14519 11339
rect 14461 11299 14519 11305
rect 9401 11271 9459 11277
rect 9401 11237 9413 11271
rect 9447 11268 9459 11271
rect 10413 11271 10471 11277
rect 9447 11240 9812 11268
rect 9447 11237 9459 11240
rect 9401 11231 9459 11237
rect 6178 11160 6184 11212
rect 6236 11160 6242 11212
rect 6457 11203 6515 11209
rect 6457 11169 6469 11203
rect 6503 11200 6515 11203
rect 6503 11172 9352 11200
rect 6503 11169 6515 11172
rect 6457 11163 6515 11169
rect 2866 11092 2872 11144
rect 2924 11092 2930 11144
rect 5905 11135 5963 11141
rect 5905 11101 5917 11135
rect 5951 11132 5963 11135
rect 6086 11132 6092 11144
rect 5951 11104 6092 11132
rect 5951 11101 5963 11104
rect 5905 11095 5963 11101
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 9214 11092 9220 11144
rect 9272 11092 9278 11144
rect 7742 11064 7748 11076
rect 7682 11036 7748 11064
rect 7742 11024 7748 11036
rect 7800 11064 7806 11076
rect 8018 11064 8024 11076
rect 7800 11036 8024 11064
rect 7800 11024 7806 11036
rect 8018 11024 8024 11036
rect 8076 11024 8082 11076
rect 9324 11064 9352 11172
rect 9784 11144 9812 11240
rect 10413 11237 10425 11271
rect 10459 11237 10471 11271
rect 10413 11231 10471 11237
rect 11517 11271 11575 11277
rect 11517 11237 11529 11271
rect 11563 11237 11575 11271
rect 11517 11231 11575 11237
rect 10428 11200 10456 11231
rect 10428 11172 11376 11200
rect 9766 11092 9772 11144
rect 9824 11092 9830 11144
rect 9858 11092 9864 11144
rect 9916 11092 9922 11144
rect 11146 11141 11152 11144
rect 10229 11135 10287 11141
rect 10229 11101 10241 11135
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 11124 11135 11152 11141
rect 11124 11101 11136 11135
rect 11124 11095 11152 11101
rect 9950 11064 9956 11076
rect 9324 11036 9956 11064
rect 9950 11024 9956 11036
rect 10008 11064 10014 11076
rect 10244 11064 10272 11095
rect 11146 11092 11152 11095
rect 11204 11092 11210 11144
rect 11348 11141 11376 11172
rect 11422 11160 11428 11212
rect 11480 11200 11486 11212
rect 11532 11200 11560 11231
rect 12342 11200 12348 11212
rect 11480 11172 12348 11200
rect 11480 11160 11486 11172
rect 12342 11160 12348 11172
rect 12400 11200 12406 11212
rect 15381 11203 15439 11209
rect 15381 11200 15393 11203
rect 12400 11172 15393 11200
rect 12400 11160 12406 11172
rect 15381 11169 15393 11172
rect 15427 11169 15439 11203
rect 15381 11163 15439 11169
rect 15654 11160 15660 11212
rect 15712 11160 15718 11212
rect 17126 11160 17132 11212
rect 17184 11160 17190 11212
rect 11333 11135 11391 11141
rect 11333 11101 11345 11135
rect 11379 11101 11391 11135
rect 11333 11095 11391 11101
rect 14090 11092 14096 11144
rect 14148 11092 14154 11144
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11132 14335 11135
rect 14323 11104 15424 11132
rect 14323 11101 14335 11104
rect 14277 11095 14335 11101
rect 10008 11036 10272 11064
rect 10008 11024 10014 11036
rect 15396 11008 15424 11104
rect 15764 11036 16146 11064
rect 2406 10956 2412 11008
rect 2464 10996 2470 11008
rect 2685 10999 2743 11005
rect 2685 10996 2697 10999
rect 2464 10968 2697 10996
rect 2464 10956 2470 10968
rect 2685 10965 2697 10968
rect 2731 10965 2743 10999
rect 2685 10959 2743 10965
rect 6089 10999 6147 11005
rect 6089 10965 6101 10999
rect 6135 10996 6147 10999
rect 6362 10996 6368 11008
rect 6135 10968 6368 10996
rect 6135 10965 6147 10968
rect 6089 10959 6147 10965
rect 6362 10956 6368 10968
rect 6420 10956 6426 11008
rect 7834 10956 7840 11008
rect 7892 10996 7898 11008
rect 7929 10999 7987 11005
rect 7929 10996 7941 10999
rect 7892 10968 7941 10996
rect 7892 10956 7898 10968
rect 7929 10965 7941 10968
rect 7975 10965 7987 10999
rect 7929 10959 7987 10965
rect 15378 10956 15384 11008
rect 15436 10996 15442 11008
rect 15764 10996 15792 11036
rect 15436 10968 15792 10996
rect 15436 10956 15442 10968
rect 1104 10906 20859 10928
rect 1104 10854 5848 10906
rect 5900 10854 5912 10906
rect 5964 10854 5976 10906
rect 6028 10854 6040 10906
rect 6092 10854 6104 10906
rect 6156 10854 10747 10906
rect 10799 10854 10811 10906
rect 10863 10854 10875 10906
rect 10927 10854 10939 10906
rect 10991 10854 11003 10906
rect 11055 10854 15646 10906
rect 15698 10854 15710 10906
rect 15762 10854 15774 10906
rect 15826 10854 15838 10906
rect 15890 10854 15902 10906
rect 15954 10854 20545 10906
rect 20597 10854 20609 10906
rect 20661 10854 20673 10906
rect 20725 10854 20737 10906
rect 20789 10854 20801 10906
rect 20853 10854 20859 10906
rect 1104 10832 20859 10854
rect 3970 10752 3976 10804
rect 4028 10792 4034 10804
rect 8665 10795 8723 10801
rect 4028 10764 8616 10792
rect 4028 10752 4034 10764
rect 8018 10724 8024 10736
rect 7866 10696 8024 10724
rect 8018 10684 8024 10696
rect 8076 10684 8082 10736
rect 8588 10724 8616 10764
rect 8665 10761 8677 10795
rect 8711 10792 8723 10795
rect 9214 10792 9220 10804
rect 8711 10764 9220 10792
rect 8711 10761 8723 10764
rect 8665 10755 8723 10761
rect 9214 10752 9220 10764
rect 9272 10752 9278 10804
rect 10965 10795 11023 10801
rect 9416 10764 10364 10792
rect 9416 10724 9444 10764
rect 8588 10696 9444 10724
rect 9674 10684 9680 10736
rect 9732 10684 9738 10736
rect 2406 10616 2412 10668
rect 2464 10616 2470 10668
rect 6362 10616 6368 10668
rect 6420 10616 6426 10668
rect 7926 10616 7932 10668
rect 7984 10656 7990 10668
rect 8205 10659 8263 10665
rect 8205 10656 8217 10659
rect 7984 10628 8217 10656
rect 7984 10616 7990 10628
rect 8205 10625 8217 10628
rect 8251 10625 8263 10659
rect 8205 10619 8263 10625
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10625 8539 10659
rect 10336 10656 10364 10764
rect 10965 10761 10977 10795
rect 11011 10792 11023 10795
rect 11146 10792 11152 10804
rect 11011 10764 11152 10792
rect 11011 10761 11023 10764
rect 10965 10755 11023 10761
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 11701 10795 11759 10801
rect 11701 10792 11713 10795
rect 11296 10764 11713 10792
rect 11296 10752 11302 10764
rect 11701 10761 11713 10764
rect 11747 10792 11759 10795
rect 11790 10792 11796 10804
rect 11747 10764 11796 10792
rect 11747 10761 11759 10764
rect 11701 10755 11759 10761
rect 11790 10752 11796 10764
rect 11848 10752 11854 10804
rect 13955 10795 14013 10801
rect 13955 10761 13967 10795
rect 14001 10792 14013 10795
rect 14090 10792 14096 10804
rect 14001 10764 14096 10792
rect 14001 10761 14013 10764
rect 13955 10755 14013 10761
rect 14090 10752 14096 10764
rect 14148 10752 14154 10804
rect 17129 10795 17187 10801
rect 17129 10761 17141 10795
rect 17175 10792 17187 10795
rect 17586 10792 17592 10804
rect 17175 10764 17592 10792
rect 17175 10761 17187 10764
rect 17129 10755 17187 10761
rect 17586 10752 17592 10764
rect 17644 10752 17650 10804
rect 18509 10727 18567 10733
rect 18509 10693 18521 10727
rect 18555 10724 18567 10727
rect 18877 10727 18935 10733
rect 18877 10724 18889 10727
rect 18555 10696 18889 10724
rect 18555 10693 18567 10696
rect 18509 10687 18567 10693
rect 18877 10693 18889 10696
rect 18923 10693 18935 10727
rect 18877 10687 18935 10693
rect 19426 10684 19432 10736
rect 19484 10684 19490 10736
rect 11514 10656 11520 10668
rect 10336 10628 11520 10656
rect 8481 10619 8539 10625
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10588 6699 10591
rect 7834 10588 7840 10600
rect 6687 10560 7840 10588
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 7834 10548 7840 10560
rect 7892 10548 7898 10600
rect 8496 10588 8524 10619
rect 11514 10616 11520 10628
rect 11572 10616 11578 10668
rect 13884 10659 13942 10665
rect 13884 10625 13896 10659
rect 13930 10656 13942 10659
rect 14458 10656 14464 10668
rect 13930 10628 14464 10656
rect 13930 10625 13942 10628
rect 13884 10619 13942 10625
rect 14458 10616 14464 10628
rect 14516 10616 14522 10668
rect 17126 10616 17132 10668
rect 17184 10656 17190 10668
rect 17184 10628 17342 10656
rect 17184 10616 17190 10628
rect 8757 10591 8815 10597
rect 8757 10588 8769 10591
rect 8496 10560 8769 10588
rect 8389 10523 8447 10529
rect 8389 10489 8401 10523
rect 8435 10520 8447 10523
rect 8496 10520 8524 10560
rect 8757 10557 8769 10560
rect 8803 10557 8815 10591
rect 8757 10551 8815 10557
rect 9033 10591 9091 10597
rect 9033 10557 9045 10591
rect 9079 10588 9091 10591
rect 9122 10588 9128 10600
rect 9079 10560 9128 10588
rect 9079 10557 9091 10560
rect 9033 10551 9091 10557
rect 8435 10492 8524 10520
rect 8435 10489 8447 10492
rect 8389 10483 8447 10489
rect 2225 10455 2283 10461
rect 2225 10421 2237 10455
rect 2271 10452 2283 10455
rect 2314 10452 2320 10464
rect 2271 10424 2320 10452
rect 2271 10421 2283 10424
rect 2225 10415 2283 10421
rect 2314 10412 2320 10424
rect 2372 10412 2378 10464
rect 8110 10412 8116 10464
rect 8168 10412 8174 10464
rect 8772 10452 8800 10551
rect 9122 10548 9128 10560
rect 9180 10548 9186 10600
rect 9766 10548 9772 10600
rect 9824 10588 9830 10600
rect 10781 10591 10839 10597
rect 10781 10588 10793 10591
rect 9824 10560 10793 10588
rect 9824 10548 9830 10560
rect 10781 10557 10793 10560
rect 10827 10557 10839 10591
rect 10781 10551 10839 10557
rect 10962 10548 10968 10600
rect 11020 10588 11026 10600
rect 16390 10588 16396 10600
rect 11020 10560 16396 10588
rect 11020 10548 11026 10560
rect 16390 10548 16396 10560
rect 16448 10588 16454 10600
rect 17402 10588 17408 10600
rect 16448 10560 17408 10588
rect 16448 10548 16454 10560
rect 17402 10548 17408 10560
rect 17460 10548 17466 10600
rect 18598 10548 18604 10600
rect 18656 10548 18662 10600
rect 10597 10523 10655 10529
rect 10597 10489 10609 10523
rect 10643 10489 10655 10523
rect 10597 10483 10655 10489
rect 10042 10452 10048 10464
rect 8772 10424 10048 10452
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 10612 10452 10640 10483
rect 17218 10480 17224 10532
rect 17276 10520 17282 10532
rect 18141 10523 18199 10529
rect 18141 10520 18153 10523
rect 17276 10492 18153 10520
rect 17276 10480 17282 10492
rect 18141 10489 18153 10492
rect 18187 10489 18199 10523
rect 18141 10483 18199 10489
rect 10560 10424 10640 10452
rect 10560 10412 10566 10424
rect 11882 10412 11888 10464
rect 11940 10452 11946 10464
rect 12158 10452 12164 10464
rect 11940 10424 12164 10452
rect 11940 10412 11946 10424
rect 12158 10412 12164 10424
rect 12216 10452 12222 10464
rect 16574 10452 16580 10464
rect 12216 10424 16580 10452
rect 12216 10412 12222 10424
rect 16574 10412 16580 10424
rect 16632 10452 16638 10464
rect 17494 10452 17500 10464
rect 16632 10424 17500 10452
rect 16632 10412 16638 10424
rect 17494 10412 17500 10424
rect 17552 10412 17558 10464
rect 20346 10412 20352 10464
rect 20404 10412 20410 10464
rect 1104 10362 20700 10384
rect 1104 10310 3399 10362
rect 3451 10310 3463 10362
rect 3515 10310 3527 10362
rect 3579 10310 3591 10362
rect 3643 10310 3655 10362
rect 3707 10310 8298 10362
rect 8350 10310 8362 10362
rect 8414 10310 8426 10362
rect 8478 10310 8490 10362
rect 8542 10310 8554 10362
rect 8606 10310 13197 10362
rect 13249 10310 13261 10362
rect 13313 10310 13325 10362
rect 13377 10310 13389 10362
rect 13441 10310 13453 10362
rect 13505 10310 18096 10362
rect 18148 10310 18160 10362
rect 18212 10310 18224 10362
rect 18276 10310 18288 10362
rect 18340 10310 18352 10362
rect 18404 10310 20700 10362
rect 1104 10288 20700 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 1762 10248 1768 10260
rect 1627 10220 1768 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 1762 10208 1768 10220
rect 1820 10208 1826 10260
rect 7926 10208 7932 10260
rect 7984 10208 7990 10260
rect 9122 10208 9128 10260
rect 9180 10208 9186 10260
rect 9858 10208 9864 10260
rect 9916 10257 9922 10260
rect 9916 10251 9965 10257
rect 9916 10217 9919 10251
rect 9953 10217 9965 10251
rect 9916 10211 9965 10217
rect 9916 10208 9922 10211
rect 10042 10208 10048 10260
rect 10100 10248 10106 10260
rect 10100 10220 14412 10248
rect 10100 10208 10106 10220
rect 4249 10183 4307 10189
rect 4249 10149 4261 10183
rect 4295 10180 4307 10183
rect 4295 10152 4752 10180
rect 4295 10149 4307 10152
rect 4249 10143 4307 10149
rect 842 10004 848 10056
rect 900 10044 906 10056
rect 1397 10047 1455 10053
rect 1397 10044 1409 10047
rect 900 10016 1409 10044
rect 900 10004 906 10016
rect 1397 10013 1409 10016
rect 1443 10013 1455 10047
rect 1397 10007 1455 10013
rect 2314 10004 2320 10056
rect 2372 10004 2378 10056
rect 3970 10004 3976 10056
rect 4028 10044 4034 10056
rect 4724 10053 4752 10152
rect 13170 10140 13176 10192
rect 13228 10180 13234 10192
rect 13909 10183 13967 10189
rect 13228 10152 13860 10180
rect 13228 10140 13234 10152
rect 6270 10072 6276 10124
rect 6328 10112 6334 10124
rect 9401 10115 9459 10121
rect 9401 10112 9413 10115
rect 6328 10084 9413 10112
rect 6328 10072 6334 10084
rect 9401 10081 9413 10084
rect 9447 10081 9459 10115
rect 10226 10112 10232 10124
rect 9401 10075 9459 10081
rect 9508 10084 10232 10112
rect 4433 10047 4491 10053
rect 4433 10044 4445 10047
rect 4028 10016 4445 10044
rect 4028 10004 4034 10016
rect 4433 10013 4445 10016
rect 4479 10013 4491 10047
rect 4433 10007 4491 10013
rect 4674 10047 4752 10053
rect 4674 10013 4686 10047
rect 4720 10044 4752 10047
rect 4950 10047 5008 10053
rect 4950 10044 4962 10047
rect 4720 10016 4962 10044
rect 4720 10013 4732 10016
rect 4674 10007 4732 10013
rect 4950 10013 4962 10016
rect 4996 10044 5008 10047
rect 6288 10044 6316 10072
rect 4996 10016 6316 10044
rect 7745 10047 7803 10053
rect 4996 10013 5008 10016
rect 4950 10007 5008 10013
rect 7745 10013 7757 10047
rect 7791 10044 7803 10047
rect 7834 10044 7840 10056
rect 7791 10016 7840 10044
rect 7791 10013 7803 10016
rect 7745 10007 7803 10013
rect 7834 10004 7840 10016
rect 7892 10004 7898 10056
rect 9508 10053 9536 10084
rect 10226 10072 10232 10084
rect 10284 10112 10290 10124
rect 11057 10115 11115 10121
rect 10284 10084 10824 10112
rect 10284 10072 10290 10084
rect 9493 10047 9551 10053
rect 9493 10013 9505 10047
rect 9539 10013 9551 10047
rect 9493 10007 9551 10013
rect 10010 10047 10068 10053
rect 10010 10013 10022 10047
rect 10056 10044 10068 10047
rect 10502 10044 10508 10056
rect 10056 10016 10508 10044
rect 10056 10013 10068 10016
rect 10010 10007 10068 10013
rect 10502 10004 10508 10016
rect 10560 10004 10566 10056
rect 10796 10044 10824 10084
rect 11057 10081 11069 10115
rect 11103 10112 11115 10115
rect 11238 10112 11244 10124
rect 11103 10084 11244 10112
rect 11103 10081 11115 10084
rect 11057 10075 11115 10081
rect 11238 10072 11244 10084
rect 11296 10072 11302 10124
rect 11333 10115 11391 10121
rect 11333 10081 11345 10115
rect 11379 10112 11391 10115
rect 11701 10115 11759 10121
rect 11701 10112 11713 10115
rect 11379 10084 11713 10112
rect 11379 10081 11391 10084
rect 11333 10075 11391 10081
rect 11701 10081 11713 10084
rect 11747 10081 11759 10115
rect 11701 10075 11759 10081
rect 13078 10072 13084 10124
rect 13136 10112 13142 10124
rect 13265 10115 13323 10121
rect 13265 10112 13277 10115
rect 13136 10084 13277 10112
rect 13136 10072 13142 10084
rect 13265 10081 13277 10084
rect 13311 10081 13323 10115
rect 13265 10075 13323 10081
rect 10962 10044 10968 10056
rect 10796 10016 10968 10044
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 11422 10004 11428 10056
rect 11480 10004 11486 10056
rect 13449 10047 13507 10053
rect 13004 10016 13400 10044
rect 1949 9979 2007 9985
rect 1949 9945 1961 9979
rect 1995 9976 2007 9979
rect 2958 9976 2964 9988
rect 1995 9948 2964 9976
rect 1995 9945 2007 9948
rect 1949 9939 2007 9945
rect 2958 9936 2964 9948
rect 3016 9936 3022 9988
rect 12158 9936 12164 9988
rect 12216 9936 12222 9988
rect 4522 9868 4528 9920
rect 4580 9917 4586 9920
rect 4580 9911 4629 9917
rect 4580 9877 4583 9911
rect 4617 9877 4629 9911
rect 4580 9871 4629 9877
rect 4580 9868 4586 9871
rect 4706 9868 4712 9920
rect 4764 9908 4770 9920
rect 4847 9911 4905 9917
rect 4847 9908 4859 9911
rect 4764 9880 4859 9908
rect 4764 9868 4770 9880
rect 4847 9877 4859 9880
rect 4893 9877 4905 9911
rect 4847 9871 4905 9877
rect 11514 9868 11520 9920
rect 11572 9908 11578 9920
rect 13004 9908 13032 10016
rect 11572 9880 13032 9908
rect 13372 9908 13400 10016
rect 13449 10013 13461 10047
rect 13495 10013 13507 10047
rect 13449 10007 13507 10013
rect 13464 9976 13492 10007
rect 13538 10004 13544 10056
rect 13596 10004 13602 10056
rect 13722 10004 13728 10056
rect 13780 10004 13786 10056
rect 13832 10044 13860 10152
rect 13909 10149 13921 10183
rect 13955 10180 13967 10183
rect 14384 10180 14412 10220
rect 14458 10208 14464 10260
rect 14516 10208 14522 10260
rect 17129 10251 17187 10257
rect 17129 10217 17141 10251
rect 17175 10248 17187 10251
rect 17218 10248 17224 10260
rect 17175 10220 17224 10248
rect 17175 10217 17187 10220
rect 17129 10211 17187 10217
rect 17218 10208 17224 10220
rect 17276 10208 17282 10260
rect 13955 10152 14320 10180
rect 14384 10152 14780 10180
rect 13955 10149 13967 10152
rect 13909 10143 13967 10149
rect 14292 10121 14320 10152
rect 14752 10121 14780 10152
rect 17586 10140 17592 10192
rect 17644 10180 17650 10192
rect 18141 10183 18199 10189
rect 18141 10180 18153 10183
rect 17644 10152 18153 10180
rect 17644 10140 17650 10152
rect 18141 10149 18153 10152
rect 18187 10149 18199 10183
rect 18141 10143 18199 10149
rect 20162 10140 20168 10192
rect 20220 10140 20226 10192
rect 14093 10115 14151 10121
rect 14093 10081 14105 10115
rect 14139 10081 14151 10115
rect 14093 10075 14151 10081
rect 14277 10115 14335 10121
rect 14277 10081 14289 10115
rect 14323 10081 14335 10115
rect 14277 10075 14335 10081
rect 14737 10115 14795 10121
rect 14737 10081 14749 10115
rect 14783 10081 14795 10115
rect 14737 10075 14795 10081
rect 16485 10115 16543 10121
rect 16485 10081 16497 10115
rect 16531 10081 16543 10115
rect 16485 10075 16543 10081
rect 14108 10044 14136 10075
rect 13832 10016 14136 10044
rect 14292 9976 14320 10075
rect 16500 10044 16528 10075
rect 17402 10072 17408 10124
rect 17460 10072 17466 10124
rect 16500 10016 17342 10044
rect 20346 10004 20352 10056
rect 20404 10004 20410 10056
rect 13464 9948 14320 9976
rect 15013 9979 15071 9985
rect 15013 9945 15025 9979
rect 15059 9945 15071 9979
rect 15013 9939 15071 9945
rect 15396 9948 15502 9976
rect 15028 9908 15056 9939
rect 15396 9920 15424 9948
rect 13372 9880 15056 9908
rect 11572 9868 11578 9880
rect 15378 9868 15384 9920
rect 15436 9868 15442 9920
rect 18506 9868 18512 9920
rect 18564 9868 18570 9920
rect 1104 9818 20859 9840
rect 1104 9766 5848 9818
rect 5900 9766 5912 9818
rect 5964 9766 5976 9818
rect 6028 9766 6040 9818
rect 6092 9766 6104 9818
rect 6156 9766 10747 9818
rect 10799 9766 10811 9818
rect 10863 9766 10875 9818
rect 10927 9766 10939 9818
rect 10991 9766 11003 9818
rect 11055 9766 15646 9818
rect 15698 9766 15710 9818
rect 15762 9766 15774 9818
rect 15826 9766 15838 9818
rect 15890 9766 15902 9818
rect 15954 9766 20545 9818
rect 20597 9766 20609 9818
rect 20661 9766 20673 9818
rect 20725 9766 20737 9818
rect 20789 9766 20801 9818
rect 20853 9766 20859 9818
rect 1104 9744 20859 9766
rect 9306 9664 9312 9716
rect 9364 9704 9370 9716
rect 13078 9704 13084 9716
rect 9364 9676 13084 9704
rect 9364 9664 9370 9676
rect 13078 9664 13084 9676
rect 13136 9664 13142 9716
rect 13311 9707 13369 9713
rect 13311 9673 13323 9707
rect 13357 9704 13369 9707
rect 13538 9704 13544 9716
rect 13357 9676 13544 9704
rect 13357 9673 13369 9676
rect 13311 9667 13369 9673
rect 13538 9664 13544 9676
rect 13596 9664 13602 9716
rect 4706 9596 4712 9648
rect 4764 9596 4770 9648
rect 5718 9596 5724 9648
rect 5776 9596 5782 9648
rect 2958 9528 2964 9580
rect 3016 9528 3022 9580
rect 12342 9528 12348 9580
rect 12400 9568 12406 9580
rect 12437 9571 12495 9577
rect 12437 9568 12449 9571
rect 12400 9540 12449 9568
rect 12400 9528 12406 9540
rect 12437 9537 12449 9540
rect 12483 9537 12495 9571
rect 12437 9531 12495 9537
rect 13170 9528 13176 9580
rect 13228 9577 13234 9580
rect 13228 9571 13266 9577
rect 13254 9537 13266 9571
rect 13228 9531 13266 9537
rect 13228 9528 13234 9531
rect 1670 9460 1676 9512
rect 1728 9460 1734 9512
rect 3878 9460 3884 9512
rect 3936 9500 3942 9512
rect 4433 9503 4491 9509
rect 4433 9500 4445 9503
rect 3936 9472 4445 9500
rect 3936 9460 3942 9472
rect 4433 9469 4445 9472
rect 4479 9500 4491 9503
rect 6181 9503 6239 9509
rect 4479 9472 5764 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 5736 9432 5764 9472
rect 6181 9469 6193 9503
rect 6227 9500 6239 9503
rect 7190 9500 7196 9512
rect 6227 9472 7196 9500
rect 6227 9469 6239 9472
rect 6181 9463 6239 9469
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 6638 9432 6644 9444
rect 5736 9404 6644 9432
rect 6638 9392 6644 9404
rect 6696 9392 6702 9444
rect 12621 9435 12679 9441
rect 12621 9401 12633 9435
rect 12667 9432 12679 9435
rect 13722 9432 13728 9444
rect 12667 9404 13728 9432
rect 12667 9401 12679 9404
rect 12621 9395 12679 9401
rect 13722 9392 13728 9404
rect 13780 9392 13786 9444
rect 1104 9274 20700 9296
rect 1104 9222 3399 9274
rect 3451 9222 3463 9274
rect 3515 9222 3527 9274
rect 3579 9222 3591 9274
rect 3643 9222 3655 9274
rect 3707 9222 8298 9274
rect 8350 9222 8362 9274
rect 8414 9222 8426 9274
rect 8478 9222 8490 9274
rect 8542 9222 8554 9274
rect 8606 9222 13197 9274
rect 13249 9222 13261 9274
rect 13313 9222 13325 9274
rect 13377 9222 13389 9274
rect 13441 9222 13453 9274
rect 13505 9222 18096 9274
rect 18148 9222 18160 9274
rect 18212 9222 18224 9274
rect 18276 9222 18288 9274
rect 18340 9222 18352 9274
rect 18404 9222 20700 9274
rect 1104 9200 20700 9222
rect 5626 9120 5632 9172
rect 5684 9120 5690 9172
rect 3878 8984 3884 9036
rect 3936 8984 3942 9036
rect 4157 9027 4215 9033
rect 4157 8993 4169 9027
rect 4203 9024 4215 9027
rect 4522 9024 4528 9036
rect 4203 8996 4528 9024
rect 4203 8993 4215 8996
rect 4157 8987 4215 8993
rect 4522 8984 4528 8996
rect 4580 8984 4586 9036
rect 7006 8916 7012 8968
rect 7064 8956 7070 8968
rect 7101 8959 7159 8965
rect 7101 8956 7113 8959
rect 7064 8928 7113 8956
rect 7064 8916 7070 8928
rect 7101 8925 7113 8928
rect 7147 8925 7159 8959
rect 7101 8919 7159 8925
rect 7558 8916 7564 8968
rect 7616 8956 7622 8968
rect 8110 8956 8116 8968
rect 7616 8928 8116 8956
rect 7616 8916 7622 8928
rect 8110 8916 8116 8928
rect 8168 8916 8174 8968
rect 20346 8916 20352 8968
rect 20404 8916 20410 8968
rect 4798 8848 4804 8900
rect 4856 8848 4862 8900
rect 6733 8891 6791 8897
rect 6733 8857 6745 8891
rect 6779 8888 6791 8891
rect 6779 8860 7420 8888
rect 6779 8857 6791 8860
rect 6733 8851 6791 8857
rect 6638 8780 6644 8832
rect 6696 8780 6702 8832
rect 7190 8780 7196 8832
rect 7248 8780 7254 8832
rect 7392 8829 7420 8860
rect 7377 8823 7435 8829
rect 7377 8789 7389 8823
rect 7423 8789 7435 8823
rect 7377 8783 7435 8789
rect 20162 8780 20168 8832
rect 20220 8780 20226 8832
rect 1104 8730 20859 8752
rect 1104 8678 5848 8730
rect 5900 8678 5912 8730
rect 5964 8678 5976 8730
rect 6028 8678 6040 8730
rect 6092 8678 6104 8730
rect 6156 8678 10747 8730
rect 10799 8678 10811 8730
rect 10863 8678 10875 8730
rect 10927 8678 10939 8730
rect 10991 8678 11003 8730
rect 11055 8678 15646 8730
rect 15698 8678 15710 8730
rect 15762 8678 15774 8730
rect 15826 8678 15838 8730
rect 15890 8678 15902 8730
rect 15954 8678 20545 8730
rect 20597 8678 20609 8730
rect 20661 8678 20673 8730
rect 20725 8678 20737 8730
rect 20789 8678 20801 8730
rect 20853 8678 20859 8730
rect 1104 8656 20859 8678
rect 13357 8619 13415 8625
rect 13357 8585 13369 8619
rect 13403 8585 13415 8619
rect 13357 8579 13415 8585
rect 7282 8440 7288 8492
rect 7340 8440 7346 8492
rect 9154 8466 9628 8480
rect 9140 8452 9628 8466
rect 7745 8415 7803 8421
rect 7745 8381 7757 8415
rect 7791 8381 7803 8415
rect 7745 8375 7803 8381
rect 8021 8415 8079 8421
rect 8021 8381 8033 8415
rect 8067 8412 8079 8415
rect 8662 8412 8668 8424
rect 8067 8384 8668 8412
rect 8067 8381 8079 8384
rect 8021 8375 8079 8381
rect 7469 8347 7527 8353
rect 7469 8313 7481 8347
rect 7515 8344 7527 8347
rect 7760 8344 7788 8375
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 7515 8316 7788 8344
rect 7515 8313 7527 8316
rect 7469 8307 7527 8313
rect 8018 8236 8024 8288
rect 8076 8276 8082 8288
rect 9140 8276 9168 8452
rect 8076 8248 9168 8276
rect 8076 8236 8082 8248
rect 9490 8236 9496 8288
rect 9548 8236 9554 8288
rect 9600 8276 9628 8452
rect 11882 8440 11888 8492
rect 11940 8480 11946 8492
rect 11977 8483 12035 8489
rect 11977 8480 11989 8483
rect 11940 8452 11989 8480
rect 11940 8440 11946 8452
rect 11977 8449 11989 8452
rect 12023 8449 12035 8483
rect 11977 8443 12035 8449
rect 12345 8483 12403 8489
rect 12345 8449 12357 8483
rect 12391 8480 12403 8483
rect 12434 8480 12440 8492
rect 12391 8452 12440 8480
rect 12391 8449 12403 8452
rect 12345 8443 12403 8449
rect 12434 8440 12440 8452
rect 12492 8440 12498 8492
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 13173 8483 13231 8489
rect 13173 8480 13185 8483
rect 12584 8452 13185 8480
rect 12584 8440 12590 8452
rect 13173 8449 13185 8452
rect 13219 8449 13231 8483
rect 13372 8480 13400 8579
rect 16022 8576 16028 8628
rect 16080 8616 16086 8628
rect 16206 8616 16212 8628
rect 16080 8588 16212 8616
rect 16080 8576 16086 8588
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 20346 8576 20352 8628
rect 20404 8576 20410 8628
rect 18414 8548 18420 8560
rect 16960 8520 18420 8548
rect 14093 8483 14151 8489
rect 14093 8480 14105 8483
rect 13372 8452 14105 8480
rect 13173 8443 13231 8449
rect 14093 8449 14105 8452
rect 14139 8480 14151 8483
rect 14369 8483 14427 8489
rect 14369 8480 14381 8483
rect 14139 8452 14381 8480
rect 14139 8449 14151 8452
rect 14093 8443 14151 8449
rect 14369 8449 14381 8452
rect 14415 8449 14427 8483
rect 14369 8443 14427 8449
rect 15470 8440 15476 8492
rect 15528 8480 15534 8492
rect 16960 8489 16988 8520
rect 18414 8508 18420 8520
rect 18472 8508 18478 8560
rect 18506 8508 18512 8560
rect 18564 8548 18570 8560
rect 18877 8551 18935 8557
rect 18877 8548 18889 8551
rect 18564 8520 18889 8548
rect 18564 8508 18570 8520
rect 18877 8517 18889 8520
rect 18923 8517 18935 8551
rect 18877 8511 18935 8517
rect 19426 8508 19432 8560
rect 19484 8508 19490 8560
rect 15841 8483 15899 8489
rect 15841 8480 15853 8483
rect 15528 8452 15853 8480
rect 15528 8440 15534 8452
rect 15841 8449 15853 8452
rect 15887 8449 15899 8483
rect 15841 8443 15899 8449
rect 16945 8483 17003 8489
rect 16945 8449 16957 8483
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 17218 8440 17224 8492
rect 17276 8440 17282 8492
rect 17862 8440 17868 8492
rect 17920 8440 17926 8492
rect 18049 8483 18107 8489
rect 18049 8449 18061 8483
rect 18095 8480 18107 8483
rect 18141 8483 18199 8489
rect 18141 8480 18153 8483
rect 18095 8452 18153 8480
rect 18095 8449 18107 8452
rect 18049 8443 18107 8449
rect 18141 8449 18153 8452
rect 18187 8449 18199 8483
rect 18141 8443 18199 8449
rect 17678 8372 17684 8424
rect 17736 8372 17742 8424
rect 18598 8372 18604 8424
rect 18656 8372 18662 8424
rect 14553 8347 14611 8353
rect 14553 8313 14565 8347
rect 14599 8344 14611 8347
rect 16298 8344 16304 8356
rect 14599 8316 16304 8344
rect 14599 8313 14611 8316
rect 14553 8307 14611 8313
rect 16298 8304 16304 8316
rect 16356 8304 16362 8356
rect 17129 8347 17187 8353
rect 17129 8313 17141 8347
rect 17175 8344 17187 8347
rect 17954 8344 17960 8356
rect 17175 8316 17960 8344
rect 17175 8313 17187 8316
rect 17129 8307 17187 8313
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 10502 8276 10508 8288
rect 9600 8248 10508 8276
rect 10502 8236 10508 8248
rect 10560 8236 10566 8288
rect 11790 8236 11796 8288
rect 11848 8236 11854 8288
rect 11974 8236 11980 8288
rect 12032 8276 12038 8288
rect 12161 8279 12219 8285
rect 12161 8276 12173 8279
rect 12032 8248 12173 8276
rect 12032 8236 12038 8248
rect 12161 8245 12173 8248
rect 12207 8245 12219 8279
rect 12161 8239 12219 8245
rect 14274 8236 14280 8288
rect 14332 8236 14338 8288
rect 17310 8236 17316 8288
rect 17368 8276 17374 8288
rect 17405 8279 17463 8285
rect 17405 8276 17417 8279
rect 17368 8248 17417 8276
rect 17368 8236 17374 8248
rect 17405 8245 17417 8248
rect 17451 8245 17463 8279
rect 17405 8239 17463 8245
rect 18325 8279 18383 8285
rect 18325 8245 18337 8279
rect 18371 8276 18383 8279
rect 18414 8276 18420 8288
rect 18371 8248 18420 8276
rect 18371 8245 18383 8248
rect 18325 8239 18383 8245
rect 18414 8236 18420 8248
rect 18472 8236 18478 8288
rect 1104 8186 20700 8208
rect 1104 8134 3399 8186
rect 3451 8134 3463 8186
rect 3515 8134 3527 8186
rect 3579 8134 3591 8186
rect 3643 8134 3655 8186
rect 3707 8134 8298 8186
rect 8350 8134 8362 8186
rect 8414 8134 8426 8186
rect 8478 8134 8490 8186
rect 8542 8134 8554 8186
rect 8606 8134 13197 8186
rect 13249 8134 13261 8186
rect 13313 8134 13325 8186
rect 13377 8134 13389 8186
rect 13441 8134 13453 8186
rect 13505 8134 18096 8186
rect 18148 8134 18160 8186
rect 18212 8134 18224 8186
rect 18276 8134 18288 8186
rect 18340 8134 18352 8186
rect 18404 8134 20700 8186
rect 1104 8112 20700 8134
rect 3234 8032 3240 8084
rect 3292 8032 3298 8084
rect 8389 8075 8447 8081
rect 8389 8041 8401 8075
rect 8435 8072 8447 8075
rect 8662 8072 8668 8084
rect 8435 8044 8668 8072
rect 8435 8041 8447 8044
rect 8389 8035 8447 8041
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 9030 8032 9036 8084
rect 9088 8072 9094 8084
rect 9088 8044 11744 8072
rect 9088 8032 9094 8044
rect 6270 8004 6276 8016
rect 2884 7976 6276 8004
rect 2884 7880 2912 7976
rect 6270 7964 6276 7976
rect 6328 7964 6334 8016
rect 6549 8007 6607 8013
rect 6549 7973 6561 8007
rect 6595 7973 6607 8007
rect 9401 8007 9459 8013
rect 9401 8004 9413 8007
rect 6549 7967 6607 7973
rect 8956 7976 9413 8004
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 4338 7936 4344 7948
rect 4111 7908 4344 7936
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7868 2375 7871
rect 2774 7868 2780 7880
rect 2363 7840 2780 7868
rect 2363 7837 2375 7840
rect 2317 7831 2375 7837
rect 2774 7828 2780 7840
rect 2832 7828 2838 7880
rect 2866 7828 2872 7880
rect 2924 7828 2930 7880
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7837 3019 7871
rect 2961 7831 3019 7837
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7837 3479 7871
rect 3421 7831 3479 7837
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7868 3663 7871
rect 3835 7871 3893 7877
rect 3835 7868 3847 7871
rect 3651 7840 3847 7868
rect 3651 7837 3663 7840
rect 3605 7831 3663 7837
rect 3835 7837 3847 7840
rect 3881 7837 3893 7871
rect 3835 7831 3893 7837
rect 3938 7871 3996 7877
rect 3938 7837 3950 7871
rect 3984 7868 3996 7871
rect 4080 7868 4108 7899
rect 4338 7896 4344 7908
rect 4396 7896 4402 7948
rect 6564 7936 6592 7967
rect 6641 7939 6699 7945
rect 6641 7936 6653 7939
rect 4908 7908 6500 7936
rect 6564 7908 6653 7936
rect 4908 7877 4936 7908
rect 3984 7840 4108 7868
rect 4249 7871 4307 7877
rect 3984 7837 3996 7840
rect 3938 7831 3996 7837
rect 4249 7837 4261 7871
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7837 4951 7871
rect 4893 7831 4951 7837
rect 5077 7871 5135 7877
rect 5077 7837 5089 7871
rect 5123 7868 5135 7871
rect 5215 7871 5273 7877
rect 5215 7868 5227 7871
rect 5123 7840 5227 7868
rect 5123 7837 5135 7840
rect 5077 7831 5135 7837
rect 5215 7837 5227 7840
rect 5261 7837 5273 7871
rect 5215 7831 5273 7837
rect 5318 7871 5376 7877
rect 5318 7837 5330 7871
rect 5364 7868 5376 7871
rect 6365 7871 6423 7877
rect 5364 7837 5396 7868
rect 5318 7831 5396 7837
rect 6365 7837 6377 7871
rect 6411 7837 6423 7871
rect 6365 7831 6423 7837
rect 2976 7800 3004 7831
rect 3436 7800 3464 7831
rect 4264 7800 4292 7831
rect 2516 7772 3004 7800
rect 3160 7772 4292 7800
rect 4433 7803 4491 7809
rect 2516 7741 2544 7772
rect 2501 7735 2559 7741
rect 2501 7701 2513 7735
rect 2547 7701 2559 7735
rect 2501 7695 2559 7701
rect 2590 7692 2596 7744
rect 2648 7732 2654 7744
rect 3160 7741 3188 7772
rect 4433 7769 4445 7803
rect 4479 7800 4491 7803
rect 5368 7800 5396 7831
rect 4479 7772 5396 7800
rect 4479 7769 4491 7772
rect 4433 7763 4491 7769
rect 2685 7735 2743 7741
rect 2685 7732 2697 7735
rect 2648 7704 2697 7732
rect 2648 7692 2654 7704
rect 2685 7701 2697 7704
rect 2731 7701 2743 7735
rect 2685 7695 2743 7701
rect 3145 7735 3203 7741
rect 3145 7701 3157 7735
rect 3191 7701 3203 7735
rect 3145 7695 3203 7701
rect 4709 7735 4767 7741
rect 4709 7701 4721 7735
rect 4755 7732 4767 7735
rect 4798 7732 4804 7744
rect 4755 7704 4804 7732
rect 4755 7701 4767 7704
rect 4709 7695 4767 7701
rect 4798 7692 4804 7704
rect 4856 7692 4862 7744
rect 6380 7732 6408 7831
rect 6472 7800 6500 7908
rect 6641 7905 6653 7908
rect 6687 7905 6699 7939
rect 6641 7899 6699 7905
rect 6917 7939 6975 7945
rect 6917 7905 6929 7939
rect 6963 7936 6975 7939
rect 7558 7936 7564 7948
rect 6963 7908 7564 7936
rect 6963 7905 6975 7908
rect 6917 7899 6975 7905
rect 7558 7896 7564 7908
rect 7616 7896 7622 7948
rect 8018 7828 8024 7880
rect 8076 7828 8082 7880
rect 8956 7877 8984 7976
rect 9401 7973 9413 7976
rect 9447 7973 9459 8007
rect 9401 7967 9459 7973
rect 9861 8007 9919 8013
rect 9861 7973 9873 8007
rect 9907 7973 9919 8007
rect 9861 7967 9919 7973
rect 8941 7871 8999 7877
rect 8941 7837 8953 7871
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7837 9275 7871
rect 9416 7868 9444 7967
rect 9876 7936 9904 7967
rect 10137 7939 10195 7945
rect 10137 7936 10149 7939
rect 9876 7908 10149 7936
rect 10137 7905 10149 7908
rect 10183 7905 10195 7939
rect 10137 7899 10195 7905
rect 9677 7871 9735 7877
rect 9677 7868 9689 7871
rect 9416 7840 9689 7868
rect 9217 7831 9275 7837
rect 9677 7837 9689 7840
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 6914 7800 6920 7812
rect 6472 7772 6920 7800
rect 6914 7760 6920 7772
rect 6972 7760 6978 7812
rect 8202 7760 8208 7812
rect 8260 7800 8266 7812
rect 9232 7800 9260 7831
rect 8260 7772 9260 7800
rect 8260 7760 8266 7772
rect 7282 7732 7288 7744
rect 6380 7704 7288 7732
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 9122 7692 9128 7744
rect 9180 7692 9186 7744
rect 9232 7732 9260 7772
rect 10410 7760 10416 7812
rect 10468 7760 10474 7812
rect 10502 7760 10508 7812
rect 10560 7800 10566 7812
rect 11716 7800 11744 8044
rect 11882 8032 11888 8084
rect 11940 8032 11946 8084
rect 18049 8075 18107 8081
rect 18049 8041 18061 8075
rect 18095 8072 18107 8075
rect 18506 8072 18512 8084
rect 18095 8044 18512 8072
rect 18095 8041 18107 8044
rect 18049 8035 18107 8041
rect 18506 8032 18512 8044
rect 18564 8032 18570 8084
rect 11900 8004 11928 8032
rect 16209 8007 16267 8013
rect 11900 7976 12112 8004
rect 11974 7896 11980 7948
rect 12032 7896 12038 7948
rect 12084 7936 12112 7976
rect 16209 7973 16221 8007
rect 16255 8004 16267 8007
rect 16255 7976 16436 8004
rect 16255 7973 16267 7976
rect 16209 7967 16267 7973
rect 12253 7939 12311 7945
rect 12253 7936 12265 7939
rect 12084 7908 12265 7936
rect 12253 7905 12265 7908
rect 12299 7905 12311 7939
rect 12253 7899 12311 7905
rect 14274 7896 14280 7948
rect 14332 7936 14338 7948
rect 14461 7939 14519 7945
rect 14461 7936 14473 7939
rect 14332 7908 14473 7936
rect 14332 7896 14338 7908
rect 14461 7905 14473 7908
rect 14507 7905 14519 7939
rect 14461 7899 14519 7905
rect 16298 7896 16304 7948
rect 16356 7896 16362 7948
rect 16408 7936 16436 7976
rect 16574 7936 16580 7948
rect 16408 7908 16580 7936
rect 16574 7896 16580 7908
rect 16632 7896 16638 7948
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7868 18291 7871
rect 18414 7868 18420 7880
rect 18279 7840 18420 7868
rect 18279 7837 18291 7840
rect 18233 7831 18291 7837
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 12710 7800 12716 7812
rect 10560 7772 10902 7800
rect 11716 7772 12716 7800
rect 10560 7760 10566 7772
rect 12710 7760 12716 7772
rect 12768 7760 12774 7812
rect 14734 7760 14740 7812
rect 14792 7760 14798 7812
rect 14844 7772 15226 7800
rect 16684 7772 17066 7800
rect 12526 7732 12532 7744
rect 9232 7704 12532 7732
rect 12526 7692 12532 7704
rect 12584 7692 12590 7744
rect 13725 7735 13783 7741
rect 13725 7701 13737 7735
rect 13771 7732 13783 7735
rect 13906 7732 13912 7744
rect 13771 7704 13912 7732
rect 13771 7701 13783 7704
rect 13725 7695 13783 7701
rect 13906 7692 13912 7704
rect 13964 7692 13970 7744
rect 14090 7692 14096 7744
rect 14148 7732 14154 7744
rect 14844 7732 14872 7772
rect 14148 7704 14872 7732
rect 15120 7732 15148 7772
rect 16684 7732 16712 7772
rect 18598 7760 18604 7812
rect 18656 7760 18662 7812
rect 15120 7704 16712 7732
rect 14148 7692 14154 7704
rect 1104 7642 20859 7664
rect 1104 7590 5848 7642
rect 5900 7590 5912 7642
rect 5964 7590 5976 7642
rect 6028 7590 6040 7642
rect 6092 7590 6104 7642
rect 6156 7590 10747 7642
rect 10799 7590 10811 7642
rect 10863 7590 10875 7642
rect 10927 7590 10939 7642
rect 10991 7590 11003 7642
rect 11055 7590 15646 7642
rect 15698 7590 15710 7642
rect 15762 7590 15774 7642
rect 15826 7590 15838 7642
rect 15890 7590 15902 7642
rect 15954 7590 20545 7642
rect 20597 7590 20609 7642
rect 20661 7590 20673 7642
rect 20725 7590 20737 7642
rect 20789 7590 20801 7642
rect 20853 7590 20859 7642
rect 1104 7568 20859 7590
rect 4246 7528 4252 7540
rect 2608 7500 4252 7528
rect 2608 7460 2636 7500
rect 4246 7488 4252 7500
rect 4304 7488 4310 7540
rect 4338 7488 4344 7540
rect 4396 7528 4402 7540
rect 5077 7531 5135 7537
rect 5077 7528 5089 7531
rect 4396 7500 5089 7528
rect 4396 7488 4402 7500
rect 5077 7497 5089 7500
rect 5123 7497 5135 7531
rect 5077 7491 5135 7497
rect 7193 7531 7251 7537
rect 7193 7497 7205 7531
rect 7239 7528 7251 7531
rect 7282 7528 7288 7540
rect 7239 7500 7288 7528
rect 7239 7497 7251 7500
rect 7193 7491 7251 7497
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 10410 7488 10416 7540
rect 10468 7528 10474 7540
rect 10873 7531 10931 7537
rect 10873 7528 10885 7531
rect 10468 7500 10885 7528
rect 10468 7488 10474 7500
rect 10873 7497 10885 7500
rect 10919 7497 10931 7531
rect 10873 7491 10931 7497
rect 2530 7432 2636 7460
rect 3142 7420 3148 7472
rect 3200 7460 3206 7472
rect 3605 7463 3663 7469
rect 3605 7460 3617 7463
rect 3200 7432 3617 7460
rect 3200 7420 3206 7432
rect 3605 7429 3617 7432
rect 3651 7429 3663 7463
rect 5350 7460 5356 7472
rect 4830 7432 5356 7460
rect 3605 7423 3663 7429
rect 5350 7420 5356 7432
rect 5408 7420 5414 7472
rect 9401 7463 9459 7469
rect 9401 7429 9413 7463
rect 9447 7460 9459 7463
rect 9490 7460 9496 7472
rect 9447 7432 9496 7460
rect 9447 7429 9459 7432
rect 9401 7423 9459 7429
rect 9490 7420 9496 7432
rect 9548 7420 9554 7472
rect 2774 7352 2780 7404
rect 2832 7392 2838 7404
rect 2832 7364 3004 7392
rect 2832 7352 2838 7364
rect 2866 7284 2872 7336
rect 2924 7284 2930 7336
rect 2976 7324 3004 7364
rect 3234 7352 3240 7404
rect 3292 7352 3298 7404
rect 7190 7352 7196 7404
rect 7248 7392 7254 7404
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 7248 7364 7389 7392
rect 7248 7352 7254 7364
rect 7377 7361 7389 7364
rect 7423 7392 7435 7395
rect 8202 7392 8208 7404
rect 7423 7364 8208 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 9122 7352 9128 7404
rect 9180 7352 9186 7404
rect 10502 7352 10508 7404
rect 10560 7352 10566 7404
rect 10888 7392 10916 7491
rect 12434 7488 12440 7540
rect 12492 7488 12498 7540
rect 12710 7488 12716 7540
rect 12768 7488 12774 7540
rect 14090 7528 14096 7540
rect 13832 7500 14096 7528
rect 11790 7420 11796 7472
rect 11848 7420 11854 7472
rect 11149 7395 11207 7401
rect 11149 7392 11161 7395
rect 10888 7364 11161 7392
rect 11149 7361 11161 7364
rect 11195 7361 11207 7395
rect 11149 7355 11207 7361
rect 12253 7395 12311 7401
rect 12253 7361 12265 7395
rect 12299 7361 12311 7395
rect 12452 7392 12480 7488
rect 12728 7460 12756 7488
rect 13832 7460 13860 7500
rect 14090 7488 14096 7500
rect 14148 7488 14154 7540
rect 14734 7488 14740 7540
rect 14792 7528 14798 7540
rect 14921 7531 14979 7537
rect 14921 7528 14933 7531
rect 14792 7500 14933 7528
rect 14792 7488 14798 7500
rect 14921 7497 14933 7500
rect 14967 7497 14979 7531
rect 14921 7491 14979 7497
rect 12728 7432 13938 7460
rect 12713 7395 12771 7401
rect 12713 7392 12725 7395
rect 12452 7364 12725 7392
rect 12253 7355 12311 7361
rect 12713 7361 12725 7364
rect 12759 7361 12771 7395
rect 14936 7392 14964 7491
rect 15470 7488 15476 7540
rect 15528 7488 15534 7540
rect 16853 7531 16911 7537
rect 16853 7497 16865 7531
rect 16899 7528 16911 7531
rect 17218 7528 17224 7540
rect 16899 7500 17224 7528
rect 16899 7497 16911 7500
rect 16853 7491 16911 7497
rect 17218 7488 17224 7500
rect 17276 7488 17282 7540
rect 17678 7488 17684 7540
rect 17736 7488 17742 7540
rect 15289 7395 15347 7401
rect 15289 7392 15301 7395
rect 14936 7364 15301 7392
rect 12713 7355 12771 7361
rect 15289 7361 15301 7364
rect 15335 7361 15347 7395
rect 15289 7355 15347 7361
rect 3329 7327 3387 7333
rect 3329 7324 3341 7327
rect 2976 7296 3341 7324
rect 3329 7293 3341 7296
rect 3375 7324 3387 7327
rect 12268 7324 12296 7355
rect 16574 7352 16580 7404
rect 16632 7392 16638 7404
rect 16669 7395 16727 7401
rect 16669 7392 16681 7395
rect 16632 7364 16681 7392
rect 16632 7352 16638 7364
rect 16669 7361 16681 7364
rect 16715 7361 16727 7395
rect 16669 7355 16727 7361
rect 17310 7352 17316 7404
rect 17368 7352 17374 7404
rect 17954 7352 17960 7404
rect 18012 7352 18018 7404
rect 18598 7352 18604 7404
rect 18656 7352 18662 7404
rect 12526 7324 12532 7336
rect 3375 7296 10548 7324
rect 12268 7296 12532 7324
rect 3375 7293 3387 7296
rect 3329 7287 3387 7293
rect 10520 7268 10548 7296
rect 12526 7284 12532 7296
rect 12584 7284 12590 7336
rect 13173 7327 13231 7333
rect 13173 7293 13185 7327
rect 13219 7293 13231 7327
rect 13173 7287 13231 7293
rect 13449 7327 13507 7333
rect 13449 7293 13461 7327
rect 13495 7324 13507 7327
rect 13906 7324 13912 7336
rect 13495 7296 13912 7324
rect 13495 7293 13507 7296
rect 13449 7287 13507 7293
rect 10502 7216 10508 7268
rect 10560 7216 10566 7268
rect 12897 7259 12955 7265
rect 12897 7225 12909 7259
rect 12943 7256 12955 7259
rect 13188 7256 13216 7287
rect 13906 7284 13912 7296
rect 13964 7284 13970 7336
rect 17405 7327 17463 7333
rect 17405 7293 17417 7327
rect 17451 7293 17463 7327
rect 17405 7287 17463 7293
rect 12943 7228 13216 7256
rect 17420 7256 17448 7287
rect 18414 7284 18420 7336
rect 18472 7324 18478 7336
rect 18877 7327 18935 7333
rect 18877 7324 18889 7327
rect 18472 7296 18889 7324
rect 18472 7284 18478 7296
rect 18877 7293 18889 7296
rect 18923 7293 18935 7327
rect 18877 7287 18935 7293
rect 17773 7259 17831 7265
rect 17773 7256 17785 7259
rect 17420 7228 17785 7256
rect 12943 7225 12955 7228
rect 12897 7219 12955 7225
rect 17773 7225 17785 7228
rect 17819 7225 17831 7259
rect 17773 7219 17831 7225
rect 1443 7191 1501 7197
rect 1443 7157 1455 7191
rect 1489 7188 1501 7191
rect 1946 7188 1952 7200
rect 1489 7160 1952 7188
rect 1489 7157 1501 7160
rect 1443 7151 1501 7157
rect 1946 7148 1952 7160
rect 2004 7148 2010 7200
rect 4246 7148 4252 7200
rect 4304 7188 4310 7200
rect 5350 7188 5356 7200
rect 4304 7160 5356 7188
rect 4304 7148 4310 7160
rect 5350 7148 5356 7160
rect 5408 7148 5414 7200
rect 10962 7148 10968 7200
rect 11020 7148 11026 7200
rect 11882 7148 11888 7200
rect 11940 7148 11946 7200
rect 1104 7098 20700 7120
rect 1104 7046 3399 7098
rect 3451 7046 3463 7098
rect 3515 7046 3527 7098
rect 3579 7046 3591 7098
rect 3643 7046 3655 7098
rect 3707 7046 8298 7098
rect 8350 7046 8362 7098
rect 8414 7046 8426 7098
rect 8478 7046 8490 7098
rect 8542 7046 8554 7098
rect 8606 7046 13197 7098
rect 13249 7046 13261 7098
rect 13313 7046 13325 7098
rect 13377 7046 13389 7098
rect 13441 7046 13453 7098
rect 13505 7046 18096 7098
rect 18148 7046 18160 7098
rect 18212 7046 18224 7098
rect 18276 7046 18288 7098
rect 18340 7046 18352 7098
rect 18404 7046 20700 7098
rect 1104 7024 20700 7046
rect 2869 6987 2927 6993
rect 2869 6953 2881 6987
rect 2915 6984 2927 6987
rect 3142 6984 3148 6996
rect 2915 6956 3148 6984
rect 2915 6953 2927 6956
rect 2869 6947 2927 6953
rect 3142 6944 3148 6956
rect 3200 6944 3206 6996
rect 2590 6808 2596 6860
rect 2648 6808 2654 6860
rect 4617 6851 4675 6857
rect 4617 6817 4629 6851
rect 4663 6848 4675 6851
rect 5626 6848 5632 6860
rect 4663 6820 5632 6848
rect 4663 6817 4675 6820
rect 4617 6811 4675 6817
rect 2501 6783 2559 6789
rect 2501 6749 2513 6783
rect 2547 6780 2559 6783
rect 2774 6780 2780 6792
rect 2547 6752 2780 6780
rect 2547 6749 2559 6752
rect 2501 6743 2559 6749
rect 2774 6740 2780 6752
rect 2832 6780 2838 6792
rect 4632 6780 4660 6811
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 8481 6851 8539 6857
rect 8481 6817 8493 6851
rect 8527 6848 8539 6851
rect 8754 6848 8760 6860
rect 8527 6820 8760 6848
rect 8527 6817 8539 6820
rect 8481 6811 8539 6817
rect 8754 6808 8760 6820
rect 8812 6808 8818 6860
rect 17862 6808 17868 6860
rect 17920 6848 17926 6860
rect 19426 6848 19432 6860
rect 17920 6820 19432 6848
rect 17920 6808 17926 6820
rect 19426 6808 19432 6820
rect 19484 6808 19490 6860
rect 2832 6752 4660 6780
rect 2832 6740 2838 6752
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 6733 6783 6791 6789
rect 6733 6780 6745 6783
rect 6696 6752 6745 6780
rect 6696 6740 6702 6752
rect 6733 6749 6745 6752
rect 6779 6749 6791 6783
rect 6733 6743 6791 6749
rect 8573 6783 8631 6789
rect 8573 6749 8585 6783
rect 8619 6780 8631 6783
rect 8662 6780 8668 6792
rect 8619 6752 8668 6780
rect 8619 6749 8631 6752
rect 8573 6743 8631 6749
rect 8662 6740 8668 6752
rect 8720 6740 8726 6792
rect 10962 6740 10968 6792
rect 11020 6740 11026 6792
rect 13906 6740 13912 6792
rect 13964 6780 13970 6792
rect 14369 6783 14427 6789
rect 14369 6780 14381 6783
rect 13964 6752 14381 6780
rect 13964 6740 13970 6752
rect 14369 6749 14381 6752
rect 14415 6749 14427 6783
rect 14369 6743 14427 6749
rect 20346 6740 20352 6792
rect 20404 6740 20410 6792
rect 5350 6672 5356 6724
rect 5408 6672 5414 6724
rect 6362 6672 6368 6724
rect 6420 6672 6426 6724
rect 7006 6672 7012 6724
rect 7064 6672 7070 6724
rect 7742 6672 7748 6724
rect 7800 6672 7806 6724
rect 8754 6604 8760 6656
rect 8812 6604 8818 6656
rect 10502 6604 10508 6656
rect 10560 6644 10566 6656
rect 10781 6647 10839 6653
rect 10781 6644 10793 6647
rect 10560 6616 10793 6644
rect 10560 6604 10566 6616
rect 10781 6613 10793 6616
rect 10827 6613 10839 6647
rect 10781 6607 10839 6613
rect 14553 6647 14611 6653
rect 14553 6613 14565 6647
rect 14599 6644 14611 6647
rect 15562 6644 15568 6656
rect 14599 6616 15568 6644
rect 14599 6613 14611 6616
rect 14553 6607 14611 6613
rect 15562 6604 15568 6616
rect 15620 6604 15626 6656
rect 20162 6604 20168 6656
rect 20220 6604 20226 6656
rect 1104 6554 20859 6576
rect 1104 6502 5848 6554
rect 5900 6502 5912 6554
rect 5964 6502 5976 6554
rect 6028 6502 6040 6554
rect 6092 6502 6104 6554
rect 6156 6502 10747 6554
rect 10799 6502 10811 6554
rect 10863 6502 10875 6554
rect 10927 6502 10939 6554
rect 10991 6502 11003 6554
rect 11055 6502 15646 6554
rect 15698 6502 15710 6554
rect 15762 6502 15774 6554
rect 15826 6502 15838 6554
rect 15890 6502 15902 6554
rect 15954 6502 20545 6554
rect 20597 6502 20609 6554
rect 20661 6502 20673 6554
rect 20725 6502 20737 6554
rect 20789 6502 20801 6554
rect 20853 6502 20859 6554
rect 1104 6480 20859 6502
rect 6779 6443 6837 6449
rect 6779 6409 6791 6443
rect 6825 6440 6837 6443
rect 7006 6440 7012 6452
rect 6825 6412 7012 6440
rect 6825 6409 6837 6412
rect 6779 6403 6837 6409
rect 7006 6400 7012 6412
rect 7064 6400 7070 6452
rect 11238 6400 11244 6452
rect 11296 6440 11302 6452
rect 17402 6440 17408 6452
rect 11296 6412 17408 6440
rect 11296 6400 11302 6412
rect 17402 6400 17408 6412
rect 17460 6400 17466 6452
rect 20346 6400 20352 6452
rect 20404 6400 20410 6452
rect 19426 6332 19432 6384
rect 19484 6332 19490 6384
rect 5258 6264 5264 6316
rect 5316 6304 5322 6316
rect 6362 6304 6368 6316
rect 5316 6276 6368 6304
rect 5316 6264 5322 6276
rect 6362 6264 6368 6276
rect 6420 6304 6426 6316
rect 6708 6307 6766 6313
rect 6708 6304 6720 6307
rect 6420 6276 6720 6304
rect 6420 6264 6426 6276
rect 6708 6273 6720 6276
rect 6754 6304 6766 6307
rect 8662 6304 8668 6316
rect 6754 6276 8668 6304
rect 6754 6273 6766 6276
rect 6708 6267 6766 6273
rect 8662 6264 8668 6276
rect 8720 6264 8726 6316
rect 9401 6307 9459 6313
rect 9401 6273 9413 6307
rect 9447 6304 9459 6307
rect 9490 6304 9496 6316
rect 9447 6276 9496 6304
rect 9447 6273 9459 6276
rect 9401 6267 9459 6273
rect 9490 6264 9496 6276
rect 9548 6264 9554 6316
rect 17497 6307 17555 6313
rect 17497 6273 17509 6307
rect 17543 6304 17555 6307
rect 18414 6304 18420 6316
rect 17543 6276 18420 6304
rect 17543 6273 17555 6276
rect 17497 6267 17555 6273
rect 18414 6264 18420 6276
rect 18472 6264 18478 6316
rect 18506 6264 18512 6316
rect 18564 6304 18570 6316
rect 18601 6307 18659 6313
rect 18601 6304 18613 6307
rect 18564 6276 18613 6304
rect 18564 6264 18570 6276
rect 18601 6273 18613 6276
rect 18647 6273 18659 6307
rect 18601 6267 18659 6273
rect 18874 6196 18880 6248
rect 18932 6196 18938 6248
rect 9582 6060 9588 6112
rect 9640 6060 9646 6112
rect 15378 6060 15384 6112
rect 15436 6100 15442 6112
rect 16206 6100 16212 6112
rect 15436 6072 16212 6100
rect 15436 6060 15442 6072
rect 16206 6060 16212 6072
rect 16264 6060 16270 6112
rect 17313 6103 17371 6109
rect 17313 6069 17325 6103
rect 17359 6100 17371 6103
rect 17402 6100 17408 6112
rect 17359 6072 17408 6100
rect 17359 6069 17371 6072
rect 17313 6063 17371 6069
rect 17402 6060 17408 6072
rect 17460 6100 17466 6112
rect 17770 6100 17776 6112
rect 17460 6072 17776 6100
rect 17460 6060 17466 6072
rect 17770 6060 17776 6072
rect 17828 6060 17834 6112
rect 1104 6010 20700 6032
rect 1104 5958 3399 6010
rect 3451 5958 3463 6010
rect 3515 5958 3527 6010
rect 3579 5958 3591 6010
rect 3643 5958 3655 6010
rect 3707 5958 8298 6010
rect 8350 5958 8362 6010
rect 8414 5958 8426 6010
rect 8478 5958 8490 6010
rect 8542 5958 8554 6010
rect 8606 5958 13197 6010
rect 13249 5958 13261 6010
rect 13313 5958 13325 6010
rect 13377 5958 13389 6010
rect 13441 5958 13453 6010
rect 13505 5958 18096 6010
rect 18148 5958 18160 6010
rect 18212 5958 18224 6010
rect 18276 5958 18288 6010
rect 18340 5958 18352 6010
rect 18404 5958 20700 6010
rect 1104 5936 20700 5958
rect 10965 5899 11023 5905
rect 10965 5865 10977 5899
rect 11011 5896 11023 5899
rect 15473 5899 15531 5905
rect 11011 5868 14320 5896
rect 11011 5865 11023 5868
rect 10965 5859 11023 5865
rect 2590 5788 2596 5840
rect 2648 5828 2654 5840
rect 5258 5828 5264 5840
rect 2648 5800 5264 5828
rect 2648 5788 2654 5800
rect 2884 5769 2912 5800
rect 5258 5788 5264 5800
rect 5316 5788 5322 5840
rect 8573 5831 8631 5837
rect 8573 5797 8585 5831
rect 8619 5797 8631 5831
rect 8573 5791 8631 5797
rect 2869 5763 2927 5769
rect 2869 5729 2881 5763
rect 2915 5729 2927 5763
rect 2869 5723 2927 5729
rect 3142 5720 3148 5772
rect 3200 5720 3206 5772
rect 7006 5720 7012 5772
rect 7064 5760 7070 5772
rect 8588 5760 8616 5791
rect 8662 5788 8668 5840
rect 8720 5828 8726 5840
rect 8720 5800 9352 5828
rect 8720 5788 8726 5800
rect 9217 5763 9275 5769
rect 9217 5760 9229 5763
rect 7064 5732 9229 5760
rect 7064 5720 7070 5732
rect 9217 5729 9229 5732
rect 9263 5729 9275 5763
rect 9324 5760 9352 5800
rect 9493 5763 9551 5769
rect 9493 5760 9505 5763
rect 9324 5732 9505 5760
rect 9217 5723 9275 5729
rect 9493 5729 9505 5732
rect 9539 5729 9551 5763
rect 9493 5723 9551 5729
rect 10502 5720 10508 5772
rect 10560 5760 10566 5772
rect 10560 5732 10916 5760
rect 10560 5720 10566 5732
rect 2774 5652 2780 5704
rect 2832 5652 2838 5704
rect 4430 5652 4436 5704
rect 4488 5692 4494 5704
rect 5166 5701 5172 5704
rect 4709 5695 4767 5701
rect 4709 5692 4721 5695
rect 4488 5664 4721 5692
rect 4488 5652 4494 5664
rect 4709 5661 4721 5664
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5692 4951 5695
rect 5031 5695 5089 5701
rect 5031 5692 5043 5695
rect 4939 5664 5043 5692
rect 4939 5661 4951 5664
rect 4893 5655 4951 5661
rect 5031 5661 5043 5664
rect 5077 5661 5089 5695
rect 5031 5655 5089 5661
rect 5134 5695 5172 5701
rect 5134 5661 5146 5695
rect 5134 5655 5172 5661
rect 5166 5652 5172 5655
rect 5224 5652 5230 5704
rect 8754 5652 8760 5704
rect 8812 5652 8818 5704
rect 9766 5584 9772 5636
rect 9824 5624 9830 5636
rect 10888 5624 10916 5732
rect 11330 5720 11336 5772
rect 11388 5760 11394 5772
rect 11701 5763 11759 5769
rect 11701 5760 11713 5763
rect 11388 5732 11713 5760
rect 11388 5720 11394 5732
rect 11701 5729 11713 5732
rect 11747 5729 11759 5763
rect 11701 5723 11759 5729
rect 11238 5652 11244 5704
rect 11296 5652 11302 5704
rect 11425 5695 11483 5701
rect 11425 5661 11437 5695
rect 11471 5661 11483 5695
rect 14292 5678 14320 5868
rect 15473 5865 15485 5899
rect 15519 5896 15531 5899
rect 18874 5896 18880 5908
rect 15519 5868 18880 5896
rect 15519 5865 15531 5868
rect 15473 5859 15531 5865
rect 18874 5856 18880 5868
rect 18932 5856 18938 5908
rect 14458 5788 14464 5840
rect 14516 5828 14522 5840
rect 15105 5831 15163 5837
rect 15105 5828 15117 5831
rect 14516 5800 15117 5828
rect 14516 5788 14522 5800
rect 15105 5797 15117 5800
rect 15151 5797 15163 5831
rect 15105 5791 15163 5797
rect 15749 5831 15807 5837
rect 15749 5797 15761 5831
rect 15795 5828 15807 5831
rect 15795 5800 15884 5828
rect 15795 5797 15807 5800
rect 15749 5791 15807 5797
rect 14366 5720 14372 5772
rect 14424 5720 14430 5772
rect 15470 5720 15476 5772
rect 15528 5760 15534 5772
rect 15856 5769 15884 5800
rect 15841 5763 15899 5769
rect 15528 5732 15700 5760
rect 15528 5720 15534 5732
rect 11425 5655 11483 5661
rect 11440 5624 11468 5655
rect 15562 5652 15568 5704
rect 15620 5652 15626 5704
rect 9824 5596 9982 5624
rect 10888 5596 11468 5624
rect 9824 5584 9830 5596
rect 1394 5516 1400 5568
rect 1452 5556 1458 5568
rect 4525 5559 4583 5565
rect 4525 5556 4537 5559
rect 1452 5528 4537 5556
rect 1452 5516 1458 5528
rect 4525 5525 4537 5528
rect 4571 5525 4583 5559
rect 9876 5556 9904 5596
rect 12158 5584 12164 5636
rect 12216 5584 12222 5636
rect 15672 5624 15700 5732
rect 15841 5729 15853 5763
rect 15887 5729 15899 5763
rect 15841 5723 15899 5729
rect 16206 5720 16212 5772
rect 16264 5760 16270 5772
rect 18049 5763 18107 5769
rect 18049 5760 18061 5763
rect 16264 5732 18061 5760
rect 16264 5720 16270 5732
rect 18049 5729 18061 5732
rect 18095 5729 18107 5763
rect 18049 5723 18107 5729
rect 17770 5652 17776 5704
rect 17828 5652 17834 5704
rect 18414 5652 18420 5704
rect 18472 5692 18478 5704
rect 20073 5695 20131 5701
rect 20073 5692 20085 5695
rect 18472 5664 20085 5692
rect 18472 5652 18478 5664
rect 20073 5661 20085 5664
rect 20119 5661 20131 5695
rect 20073 5655 20131 5661
rect 16117 5627 16175 5633
rect 16117 5624 16129 5627
rect 15396 5596 15608 5624
rect 15672 5596 16129 5624
rect 11149 5559 11207 5565
rect 11149 5556 11161 5559
rect 9876 5528 11161 5556
rect 4525 5519 4583 5525
rect 11149 5525 11161 5528
rect 11195 5525 11207 5559
rect 11149 5519 11207 5525
rect 13173 5559 13231 5565
rect 13173 5525 13185 5559
rect 13219 5556 13231 5559
rect 13814 5556 13820 5568
rect 13219 5528 13820 5556
rect 13219 5525 13231 5528
rect 13173 5519 13231 5525
rect 13814 5516 13820 5528
rect 13872 5516 13878 5568
rect 14093 5559 14151 5565
rect 14093 5525 14105 5559
rect 14139 5556 14151 5559
rect 15396 5556 15424 5596
rect 14139 5528 15424 5556
rect 15580 5556 15608 5596
rect 16117 5593 16129 5596
rect 16163 5593 16175 5627
rect 16117 5587 16175 5593
rect 16206 5584 16212 5636
rect 16264 5624 16270 5636
rect 17678 5624 17684 5636
rect 16264 5596 16606 5624
rect 17420 5596 17684 5624
rect 16264 5584 16270 5596
rect 17420 5556 17448 5596
rect 17678 5584 17684 5596
rect 17736 5584 17742 5636
rect 15580 5528 17448 5556
rect 14139 5525 14151 5528
rect 14093 5519 14151 5525
rect 17586 5516 17592 5568
rect 17644 5516 17650 5568
rect 20254 5516 20260 5568
rect 20312 5516 20318 5568
rect 1104 5466 20859 5488
rect 1104 5414 5848 5466
rect 5900 5414 5912 5466
rect 5964 5414 5976 5466
rect 6028 5414 6040 5466
rect 6092 5414 6104 5466
rect 6156 5414 10747 5466
rect 10799 5414 10811 5466
rect 10863 5414 10875 5466
rect 10927 5414 10939 5466
rect 10991 5414 11003 5466
rect 11055 5414 15646 5466
rect 15698 5414 15710 5466
rect 15762 5414 15774 5466
rect 15826 5414 15838 5466
rect 15890 5414 15902 5466
rect 15954 5414 20545 5466
rect 20597 5414 20609 5466
rect 20661 5414 20673 5466
rect 20725 5414 20737 5466
rect 20789 5414 20801 5466
rect 20853 5414 20859 5466
rect 1104 5392 20859 5414
rect 5077 5355 5135 5361
rect 3068 5324 3740 5352
rect 3068 5284 3096 5324
rect 2806 5256 3096 5284
rect 3142 5244 3148 5296
rect 3200 5284 3206 5296
rect 3605 5287 3663 5293
rect 3605 5284 3617 5287
rect 3200 5256 3617 5284
rect 3200 5244 3206 5256
rect 3605 5253 3617 5256
rect 3651 5253 3663 5287
rect 3712 5284 3740 5324
rect 5077 5321 5089 5355
rect 5123 5352 5135 5355
rect 5166 5352 5172 5364
rect 5123 5324 5172 5352
rect 5123 5321 5135 5324
rect 5077 5315 5135 5321
rect 5166 5312 5172 5324
rect 5224 5312 5230 5364
rect 5537 5355 5595 5361
rect 5537 5321 5549 5355
rect 5583 5352 5595 5355
rect 5718 5352 5724 5364
rect 5583 5324 5724 5352
rect 5583 5321 5595 5324
rect 5537 5315 5595 5321
rect 5718 5312 5724 5324
rect 5776 5312 5782 5364
rect 13633 5355 13691 5361
rect 5828 5324 8800 5352
rect 4062 5284 4068 5296
rect 3712 5256 4068 5284
rect 3605 5247 3663 5253
rect 4062 5244 4068 5256
rect 4120 5244 4126 5296
rect 5626 5244 5632 5296
rect 5684 5284 5690 5296
rect 5828 5284 5856 5324
rect 7006 5284 7012 5296
rect 5684 5256 5856 5284
rect 5684 5244 5690 5256
rect 1394 5176 1400 5228
rect 1452 5176 1458 5228
rect 5353 5219 5411 5225
rect 5353 5216 5365 5219
rect 4738 5202 5365 5216
rect 4724 5188 5365 5202
rect 1765 5151 1823 5157
rect 1765 5117 1777 5151
rect 1811 5148 1823 5151
rect 2590 5148 2596 5160
rect 1811 5120 2596 5148
rect 1811 5117 1823 5120
rect 1765 5111 1823 5117
rect 2590 5108 2596 5120
rect 2648 5108 2654 5160
rect 3329 5151 3387 5157
rect 3329 5117 3341 5151
rect 3375 5117 3387 5151
rect 3329 5111 3387 5117
rect 3234 5021 3240 5024
rect 3191 5015 3240 5021
rect 3191 4981 3203 5015
rect 3237 4981 3240 5015
rect 3191 4975 3240 4981
rect 3234 4972 3240 4975
rect 3292 4972 3298 5024
rect 3344 5012 3372 5111
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 4724 5148 4752 5188
rect 5353 5185 5365 5188
rect 5399 5216 5411 5219
rect 5442 5216 5448 5228
rect 5399 5188 5448 5216
rect 5399 5185 5411 5188
rect 5353 5179 5411 5185
rect 5442 5176 5448 5188
rect 5500 5176 5506 5228
rect 5828 5225 5856 5256
rect 6472 5256 7012 5284
rect 6472 5225 6500 5256
rect 7006 5244 7012 5256
rect 7064 5244 7070 5296
rect 8662 5284 8668 5296
rect 7958 5256 8668 5284
rect 8662 5244 8668 5256
rect 8720 5244 8726 5296
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 6457 5219 6515 5225
rect 6457 5185 6469 5219
rect 6503 5185 6515 5219
rect 6457 5179 6515 5185
rect 4120 5120 4752 5148
rect 4120 5108 4126 5120
rect 5166 5108 5172 5160
rect 5224 5108 5230 5160
rect 5905 5151 5963 5157
rect 5905 5117 5917 5151
rect 5951 5148 5963 5151
rect 6270 5148 6276 5160
rect 5951 5120 6276 5148
rect 5951 5117 5963 5120
rect 5905 5111 5963 5117
rect 6270 5108 6276 5120
rect 6328 5108 6334 5160
rect 6733 5151 6791 5157
rect 6733 5148 6745 5151
rect 6564 5120 6745 5148
rect 6181 5083 6239 5089
rect 6181 5049 6193 5083
rect 6227 5080 6239 5083
rect 6564 5080 6592 5120
rect 6733 5117 6745 5120
rect 6779 5117 6791 5151
rect 8772 5148 8800 5324
rect 13633 5321 13645 5355
rect 13679 5352 13691 5355
rect 14458 5352 14464 5364
rect 13679 5324 14464 5352
rect 13679 5321 13691 5324
rect 13633 5315 13691 5321
rect 14458 5312 14464 5324
rect 14516 5312 14522 5364
rect 15013 5355 15071 5361
rect 15013 5321 15025 5355
rect 15059 5352 15071 5355
rect 15059 5324 16574 5352
rect 15059 5321 15071 5324
rect 15013 5315 15071 5321
rect 16022 5244 16028 5296
rect 16080 5284 16086 5296
rect 16301 5287 16359 5293
rect 16301 5284 16313 5287
rect 16080 5256 16313 5284
rect 16080 5244 16086 5256
rect 16301 5253 16313 5256
rect 16347 5253 16359 5287
rect 16546 5284 16574 5324
rect 18414 5312 18420 5364
rect 18472 5312 18478 5364
rect 16945 5287 17003 5293
rect 16945 5284 16957 5287
rect 16546 5256 16957 5284
rect 16301 5247 16359 5253
rect 16945 5253 16957 5256
rect 16991 5253 17003 5287
rect 19242 5284 19248 5296
rect 18170 5256 19248 5284
rect 16945 5247 17003 5253
rect 19242 5244 19248 5256
rect 19300 5244 19306 5296
rect 19334 5244 19340 5296
rect 19392 5244 19398 5296
rect 9582 5176 9588 5228
rect 9640 5176 9646 5228
rect 12250 5176 12256 5228
rect 12308 5216 12314 5228
rect 12308 5188 13846 5216
rect 12308 5176 12314 5188
rect 18506 5176 18512 5228
rect 18564 5176 18570 5228
rect 16485 5151 16543 5157
rect 8772 5134 13938 5148
rect 8772 5120 13952 5134
rect 6733 5111 6791 5117
rect 9769 5083 9827 5089
rect 9769 5080 9781 5083
rect 6227 5052 6592 5080
rect 7760 5052 9781 5080
rect 6227 5049 6239 5052
rect 6181 5043 6239 5049
rect 3786 5012 3792 5024
rect 3344 4984 3792 5012
rect 3786 4972 3792 4984
rect 3844 5012 3850 5024
rect 7760 5012 7788 5052
rect 9769 5049 9781 5052
rect 9815 5080 9827 5083
rect 10502 5080 10508 5092
rect 9815 5052 10508 5080
rect 9815 5049 9827 5052
rect 9769 5043 9827 5049
rect 10502 5040 10508 5052
rect 10560 5040 10566 5092
rect 3844 4984 7788 5012
rect 3844 4972 3850 4984
rect 8202 4972 8208 5024
rect 8260 4972 8266 5024
rect 13924 5012 13952 5120
rect 16485 5117 16497 5151
rect 16531 5148 16543 5151
rect 16669 5151 16727 5157
rect 16669 5148 16681 5151
rect 16531 5120 16681 5148
rect 16531 5117 16543 5120
rect 16485 5111 16543 5117
rect 16669 5117 16681 5120
rect 16715 5148 16727 5151
rect 18524 5148 18552 5176
rect 16715 5120 18552 5148
rect 16715 5117 16727 5120
rect 16669 5111 16727 5117
rect 18782 5108 18788 5160
rect 18840 5108 18846 5160
rect 14090 5040 14096 5092
rect 14148 5080 14154 5092
rect 14645 5083 14703 5089
rect 14645 5080 14657 5083
rect 14148 5052 14657 5080
rect 14148 5040 14154 5052
rect 14645 5049 14657 5052
rect 14691 5049 14703 5083
rect 14645 5043 14703 5049
rect 14366 5012 14372 5024
rect 13924 4984 14372 5012
rect 14366 4972 14372 4984
rect 14424 4972 14430 5024
rect 20070 4972 20076 5024
rect 20128 5012 20134 5024
rect 20257 5015 20315 5021
rect 20257 5012 20269 5015
rect 20128 4984 20269 5012
rect 20128 4972 20134 4984
rect 20257 4981 20269 4984
rect 20303 4981 20315 5015
rect 20257 4975 20315 4981
rect 1104 4922 20700 4944
rect 1104 4870 3399 4922
rect 3451 4870 3463 4922
rect 3515 4870 3527 4922
rect 3579 4870 3591 4922
rect 3643 4870 3655 4922
rect 3707 4870 8298 4922
rect 8350 4870 8362 4922
rect 8414 4870 8426 4922
rect 8478 4870 8490 4922
rect 8542 4870 8554 4922
rect 8606 4870 13197 4922
rect 13249 4870 13261 4922
rect 13313 4870 13325 4922
rect 13377 4870 13389 4922
rect 13441 4870 13453 4922
rect 13505 4870 18096 4922
rect 18148 4870 18160 4922
rect 18212 4870 18224 4922
rect 18276 4870 18288 4922
rect 18340 4870 18352 4922
rect 18404 4870 20700 4922
rect 1104 4848 20700 4870
rect 4430 4768 4436 4820
rect 4488 4768 4494 4820
rect 5166 4768 5172 4820
rect 5224 4808 5230 4820
rect 5307 4811 5365 4817
rect 5307 4808 5319 4811
rect 5224 4780 5319 4808
rect 5224 4768 5230 4780
rect 5307 4777 5319 4780
rect 5353 4777 5365 4811
rect 5307 4771 5365 4777
rect 5442 4768 5448 4820
rect 5500 4808 5506 4820
rect 8662 4808 8668 4820
rect 5500 4780 8668 4808
rect 5500 4768 5506 4780
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 12250 4768 12256 4820
rect 12308 4768 12314 4820
rect 14090 4768 14096 4820
rect 14148 4768 14154 4820
rect 15473 4811 15531 4817
rect 15473 4777 15485 4811
rect 15519 4808 15531 4811
rect 18782 4808 18788 4820
rect 15519 4780 18788 4808
rect 15519 4777 15531 4780
rect 15473 4771 15531 4777
rect 18782 4768 18788 4780
rect 18840 4768 18846 4820
rect 3973 4743 4031 4749
rect 3973 4709 3985 4743
rect 4019 4709 4031 4743
rect 3973 4703 4031 4709
rect 3786 4564 3792 4616
rect 3844 4564 3850 4616
rect 3988 4604 4016 4703
rect 4448 4672 4476 4768
rect 4801 4743 4859 4749
rect 4801 4709 4813 4743
rect 4847 4740 4859 4743
rect 5074 4740 5080 4752
rect 4847 4712 5080 4740
rect 4847 4709 4859 4712
rect 4801 4703 4859 4709
rect 5074 4700 5080 4712
rect 5132 4700 5138 4752
rect 7101 4743 7159 4749
rect 7101 4709 7113 4743
rect 7147 4709 7159 4743
rect 7101 4703 7159 4709
rect 4985 4675 5043 4681
rect 4985 4672 4997 4675
rect 4448 4644 4997 4672
rect 4985 4641 4997 4644
rect 5031 4641 5043 4675
rect 4985 4635 5043 4641
rect 4249 4607 4307 4613
rect 4249 4604 4261 4607
rect 3988 4576 4261 4604
rect 4249 4573 4261 4576
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 5169 4607 5227 4613
rect 5169 4573 5181 4607
rect 5215 4604 5227 4607
rect 5378 4607 5436 4613
rect 5378 4604 5390 4607
rect 5215 4576 5390 4604
rect 5215 4573 5227 4576
rect 5169 4567 5227 4573
rect 5378 4573 5390 4576
rect 5424 4573 5436 4607
rect 5378 4567 5436 4573
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4604 6975 4607
rect 7006 4604 7012 4616
rect 6963 4576 7012 4604
rect 6963 4573 6975 4576
rect 6917 4567 6975 4573
rect 7006 4564 7012 4576
rect 7064 4564 7070 4616
rect 7116 4604 7144 4703
rect 8202 4700 8208 4752
rect 8260 4700 8266 4752
rect 15102 4700 15108 4752
rect 15160 4700 15166 4752
rect 7745 4675 7803 4681
rect 7745 4672 7757 4675
rect 7576 4644 7757 4672
rect 7469 4607 7527 4613
rect 7469 4604 7481 4607
rect 7116 4576 7481 4604
rect 7469 4573 7481 4576
rect 7515 4573 7527 4607
rect 7469 4567 7527 4573
rect 3050 4496 3056 4548
rect 3108 4536 3114 4548
rect 7576 4536 7604 4644
rect 7745 4641 7757 4644
rect 7791 4641 7803 4675
rect 8220 4672 8248 4700
rect 8220 4644 8432 4672
rect 7745 4635 7803 4641
rect 7926 4604 7932 4616
rect 3108 4508 7604 4536
rect 7668 4576 7932 4604
rect 3108 4496 3114 4508
rect 7668 4477 7696 4576
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 8404 4613 8432 4644
rect 10502 4632 10508 4684
rect 10560 4632 10566 4684
rect 10781 4675 10839 4681
rect 10781 4641 10793 4675
rect 10827 4672 10839 4675
rect 11330 4672 11336 4684
rect 10827 4644 11336 4672
rect 10827 4641 10839 4644
rect 10781 4635 10839 4641
rect 11330 4632 11336 4644
rect 11388 4632 11394 4684
rect 14366 4632 14372 4684
rect 14424 4632 14430 4684
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4604 8171 4607
rect 8251 4607 8309 4613
rect 8251 4604 8263 4607
rect 8159 4576 8263 4604
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 8251 4573 8263 4576
rect 8297 4573 8309 4607
rect 8251 4567 8309 4573
rect 8354 4607 8432 4613
rect 8354 4573 8366 4607
rect 8400 4576 8432 4607
rect 8400 4573 8412 4576
rect 8354 4567 8412 4573
rect 13814 4564 13820 4616
rect 13872 4604 13878 4616
rect 13872 4576 14306 4604
rect 13872 4564 13878 4576
rect 12158 4536 12164 4548
rect 12006 4508 12164 4536
rect 12158 4496 12164 4508
rect 12216 4496 12222 4548
rect 7653 4471 7711 4477
rect 7653 4437 7665 4471
rect 7699 4437 7711 4471
rect 7653 4431 7711 4437
rect 1104 4378 20859 4400
rect 1104 4326 5848 4378
rect 5900 4326 5912 4378
rect 5964 4326 5976 4378
rect 6028 4326 6040 4378
rect 6092 4326 6104 4378
rect 6156 4326 10747 4378
rect 10799 4326 10811 4378
rect 10863 4326 10875 4378
rect 10927 4326 10939 4378
rect 10991 4326 11003 4378
rect 11055 4326 15646 4378
rect 15698 4326 15710 4378
rect 15762 4326 15774 4378
rect 15826 4326 15838 4378
rect 15890 4326 15902 4378
rect 15954 4326 20545 4378
rect 20597 4326 20609 4378
rect 20661 4326 20673 4378
rect 20725 4326 20737 4378
rect 20789 4326 20801 4378
rect 20853 4326 20859 4378
rect 1104 4304 20859 4326
rect 19334 4156 19340 4208
rect 19392 4156 19398 4208
rect 7926 4088 7932 4140
rect 7984 4128 7990 4140
rect 8113 4131 8171 4137
rect 8113 4128 8125 4131
rect 7984 4100 8125 4128
rect 7984 4088 7990 4100
rect 8113 4097 8125 4100
rect 8159 4097 8171 4131
rect 8113 4091 8171 4097
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4128 8355 4131
rect 8506 4131 8564 4137
rect 8506 4128 8518 4131
rect 8343 4100 8518 4128
rect 8343 4097 8355 4100
rect 8297 4091 8355 4097
rect 8506 4097 8518 4100
rect 8552 4097 8564 4131
rect 8506 4091 8564 4097
rect 18506 4088 18512 4140
rect 18564 4128 18570 4140
rect 18601 4131 18659 4137
rect 18601 4128 18613 4131
rect 18564 4100 18613 4128
rect 18564 4088 18570 4100
rect 18601 4097 18613 4100
rect 18647 4097 18659 4131
rect 18601 4091 18659 4097
rect 8202 4060 8208 4072
rect 7944 4032 8208 4060
rect 7944 4001 7972 4032
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 18877 4063 18935 4069
rect 18877 4060 18889 4063
rect 18708 4032 18889 4060
rect 7929 3995 7987 4001
rect 7929 3961 7941 3995
rect 7975 3961 7987 3995
rect 11882 3992 11888 4004
rect 7929 3955 7987 3961
rect 8128 3964 11888 3992
rect 2958 3884 2964 3936
rect 3016 3924 3022 3936
rect 3142 3924 3148 3936
rect 3016 3896 3148 3924
rect 3016 3884 3022 3896
rect 3142 3884 3148 3896
rect 3200 3924 3206 3936
rect 8128 3924 8156 3964
rect 11882 3952 11888 3964
rect 11940 3952 11946 4004
rect 17586 3952 17592 4004
rect 17644 3992 17650 4004
rect 18708 3992 18736 4032
rect 18877 4029 18889 4032
rect 18923 4029 18935 4063
rect 18877 4023 18935 4029
rect 17644 3964 18736 3992
rect 17644 3952 17650 3964
rect 3200 3896 8156 3924
rect 3200 3884 3206 3896
rect 8202 3884 8208 3936
rect 8260 3924 8266 3936
rect 8435 3927 8493 3933
rect 8435 3924 8447 3927
rect 8260 3896 8447 3924
rect 8260 3884 8266 3896
rect 8435 3893 8447 3896
rect 8481 3893 8493 3927
rect 8435 3887 8493 3893
rect 20346 3884 20352 3936
rect 20404 3884 20410 3936
rect 1104 3834 20700 3856
rect 1104 3782 3399 3834
rect 3451 3782 3463 3834
rect 3515 3782 3527 3834
rect 3579 3782 3591 3834
rect 3643 3782 3655 3834
rect 3707 3782 8298 3834
rect 8350 3782 8362 3834
rect 8414 3782 8426 3834
rect 8478 3782 8490 3834
rect 8542 3782 8554 3834
rect 8606 3782 13197 3834
rect 13249 3782 13261 3834
rect 13313 3782 13325 3834
rect 13377 3782 13389 3834
rect 13441 3782 13453 3834
rect 13505 3782 18096 3834
rect 18148 3782 18160 3834
rect 18212 3782 18224 3834
rect 18276 3782 18288 3834
rect 18340 3782 18352 3834
rect 18404 3782 20700 3834
rect 1104 3760 20700 3782
rect 7742 3680 7748 3732
rect 7800 3720 7806 3732
rect 7837 3723 7895 3729
rect 7837 3720 7849 3723
rect 7800 3692 7849 3720
rect 7800 3680 7806 3692
rect 7837 3689 7849 3692
rect 7883 3689 7895 3723
rect 7837 3683 7895 3689
rect 20254 3612 20260 3664
rect 20312 3612 20318 3664
rect 2869 3587 2927 3593
rect 2869 3553 2881 3587
rect 2915 3584 2927 3587
rect 5258 3584 5264 3596
rect 2915 3556 5264 3584
rect 2915 3553 2927 3556
rect 2869 3547 2927 3553
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 8202 3544 8208 3596
rect 8260 3544 8266 3596
rect 9784 3556 10548 3584
rect 9784 3528 9812 3556
rect 10520 3528 10548 3556
rect 10594 3544 10600 3596
rect 10652 3584 10658 3596
rect 10689 3587 10747 3593
rect 10689 3584 10701 3587
rect 10652 3556 10701 3584
rect 10652 3544 10658 3556
rect 10689 3553 10701 3556
rect 10735 3553 10747 3587
rect 10689 3547 10747 3553
rect 11057 3587 11115 3593
rect 11057 3553 11069 3587
rect 11103 3584 11115 3587
rect 11330 3584 11336 3596
rect 11103 3556 11336 3584
rect 11103 3553 11115 3556
rect 11057 3547 11115 3553
rect 11330 3544 11336 3556
rect 11388 3544 11394 3596
rect 15286 3544 15292 3596
rect 15344 3584 15350 3596
rect 15473 3587 15531 3593
rect 15473 3584 15485 3587
rect 15344 3556 15485 3584
rect 15344 3544 15350 3556
rect 15473 3553 15485 3556
rect 15519 3553 15531 3587
rect 15473 3547 15531 3553
rect 15654 3544 15660 3596
rect 15712 3584 15718 3596
rect 15841 3587 15899 3593
rect 15841 3584 15853 3587
rect 15712 3556 15853 3584
rect 15712 3544 15718 3556
rect 15841 3553 15853 3556
rect 15887 3584 15899 3587
rect 16022 3584 16028 3596
rect 15887 3556 16028 3584
rect 15887 3553 15899 3556
rect 15841 3547 15899 3553
rect 16022 3544 16028 3556
rect 16080 3544 16086 3596
rect 3142 3476 3148 3528
rect 3200 3476 3206 3528
rect 4982 3476 4988 3528
rect 5040 3476 5046 3528
rect 6914 3476 6920 3528
rect 6972 3516 6978 3528
rect 8021 3519 8079 3525
rect 8021 3516 8033 3519
rect 6972 3488 8033 3516
rect 6972 3476 6978 3488
rect 8021 3485 8033 3488
rect 8067 3516 8079 3519
rect 9766 3516 9772 3528
rect 8067 3488 9772 3516
rect 8067 3485 8079 3488
rect 8021 3479 8079 3485
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 9953 3519 10011 3525
rect 9953 3485 9965 3519
rect 9999 3516 10011 3519
rect 10318 3516 10324 3528
rect 9999 3488 10324 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 10502 3476 10508 3528
rect 10560 3476 10566 3528
rect 20070 3476 20076 3528
rect 20128 3476 20134 3528
rect 4062 3448 4068 3460
rect 2438 3420 4068 3448
rect 4062 3408 4068 3420
rect 4120 3408 4126 3460
rect 5718 3408 5724 3460
rect 5776 3408 5782 3460
rect 8662 3408 8668 3460
rect 8720 3448 8726 3460
rect 8720 3420 10272 3448
rect 8720 3408 8726 3420
rect 10244 3392 10272 3420
rect 12066 3408 12072 3460
rect 12124 3448 12130 3460
rect 16206 3448 16212 3460
rect 12124 3420 15608 3448
rect 12124 3408 12130 3420
rect 1394 3340 1400 3392
rect 1452 3340 1458 3392
rect 6733 3383 6791 3389
rect 6733 3349 6745 3383
rect 6779 3380 6791 3383
rect 7098 3380 7104 3392
rect 6779 3352 7104 3380
rect 6779 3349 6791 3352
rect 6733 3343 6791 3349
rect 7098 3340 7104 3352
rect 7156 3340 7162 3392
rect 9582 3340 9588 3392
rect 9640 3380 9646 3392
rect 9769 3383 9827 3389
rect 9769 3380 9781 3383
rect 9640 3352 9781 3380
rect 9640 3340 9646 3352
rect 9769 3349 9781 3352
rect 9815 3349 9827 3383
rect 9769 3343 9827 3349
rect 10226 3340 10232 3392
rect 10284 3340 10290 3392
rect 12526 3389 12532 3392
rect 12483 3383 12532 3389
rect 12483 3349 12495 3383
rect 12529 3349 12532 3383
rect 12483 3343 12532 3349
rect 12526 3340 12532 3343
rect 12584 3340 12590 3392
rect 15580 3380 15608 3420
rect 16132 3420 16212 3448
rect 16132 3380 16160 3420
rect 16206 3408 16212 3420
rect 16264 3408 16270 3460
rect 15580 3352 16160 3380
rect 17267 3383 17325 3389
rect 17267 3349 17279 3383
rect 17313 3380 17325 3383
rect 17402 3380 17408 3392
rect 17313 3352 17408 3380
rect 17313 3349 17325 3352
rect 17267 3343 17325 3349
rect 17402 3340 17408 3352
rect 17460 3340 17466 3392
rect 1104 3290 20859 3312
rect 1104 3238 5848 3290
rect 5900 3238 5912 3290
rect 5964 3238 5976 3290
rect 6028 3238 6040 3290
rect 6092 3238 6104 3290
rect 6156 3238 10747 3290
rect 10799 3238 10811 3290
rect 10863 3238 10875 3290
rect 10927 3238 10939 3290
rect 10991 3238 11003 3290
rect 11055 3238 15646 3290
rect 15698 3238 15710 3290
rect 15762 3238 15774 3290
rect 15826 3238 15838 3290
rect 15890 3238 15902 3290
rect 15954 3238 20545 3290
rect 20597 3238 20609 3290
rect 20661 3238 20673 3290
rect 20725 3238 20737 3290
rect 20789 3238 20801 3290
rect 20853 3238 20859 3290
rect 1104 3216 20859 3238
rect 13817 3179 13875 3185
rect 13817 3145 13829 3179
rect 13863 3176 13875 3179
rect 15102 3176 15108 3188
rect 13863 3148 15108 3176
rect 13863 3145 13875 3148
rect 13817 3139 13875 3145
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 16206 3136 16212 3188
rect 16264 3176 16270 3188
rect 16264 3148 17724 3176
rect 16264 3136 16270 3148
rect 4062 3068 4068 3120
rect 4120 3068 4126 3120
rect 7650 3068 7656 3120
rect 7708 3068 7714 3120
rect 10226 3068 10232 3120
rect 10284 3068 10290 3120
rect 12066 3068 12072 3120
rect 12124 3108 12130 3120
rect 17696 3108 17724 3148
rect 12124 3080 12834 3108
rect 17696 3080 17802 3108
rect 12124 3068 12130 3080
rect 1670 3000 1676 3052
rect 1728 3000 1734 3052
rect 4663 3043 4721 3049
rect 4663 3009 4675 3043
rect 4709 3040 4721 3043
rect 4801 3043 4859 3049
rect 4801 3040 4813 3043
rect 4709 3012 4813 3040
rect 4709 3009 4721 3012
rect 4663 3003 4721 3009
rect 4801 3009 4813 3012
rect 4847 3009 4859 3043
rect 4801 3003 4859 3009
rect 4982 3000 4988 3052
rect 5040 3040 5046 3052
rect 6638 3040 6644 3052
rect 5040 3012 6644 3040
rect 5040 3000 5046 3012
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 9306 3000 9312 3052
rect 9364 3000 9370 3052
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3040 17095 3043
rect 17126 3040 17132 3052
rect 17083 3012 17132 3040
rect 17083 3009 17095 3012
rect 17037 3003 17095 3009
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 20346 3000 20352 3052
rect 20404 3000 20410 3052
rect 2869 2975 2927 2981
rect 2869 2941 2881 2975
rect 2915 2972 2927 2975
rect 3050 2972 3056 2984
rect 2915 2944 3056 2972
rect 2915 2941 2927 2944
rect 2869 2935 2927 2941
rect 3050 2932 3056 2944
rect 3108 2932 3114 2984
rect 3237 2975 3295 2981
rect 3237 2941 3249 2975
rect 3283 2972 3295 2975
rect 5258 2972 5264 2984
rect 3283 2944 5264 2972
rect 3283 2941 3295 2944
rect 3237 2935 3295 2941
rect 5258 2932 5264 2944
rect 5316 2932 5322 2984
rect 6270 2932 6276 2984
rect 6328 2972 6334 2984
rect 6917 2975 6975 2981
rect 6917 2972 6929 2975
rect 6328 2944 6929 2972
rect 6328 2932 6334 2944
rect 6917 2941 6929 2944
rect 6963 2972 6975 2975
rect 9490 2972 9496 2984
rect 6963 2944 9496 2972
rect 6963 2941 6975 2944
rect 6917 2935 6975 2941
rect 9490 2932 9496 2944
rect 9548 2972 9554 2984
rect 9677 2975 9735 2981
rect 9677 2972 9689 2975
rect 9548 2944 9689 2972
rect 9548 2932 9554 2944
rect 9677 2941 9689 2944
rect 9723 2941 9735 2975
rect 9677 2935 9735 2941
rect 11882 2932 11888 2984
rect 11940 2972 11946 2984
rect 12069 2975 12127 2981
rect 12069 2972 12081 2975
rect 11940 2944 12081 2972
rect 11940 2932 11946 2944
rect 12069 2941 12081 2944
rect 12115 2941 12127 2975
rect 12345 2975 12403 2981
rect 12345 2972 12357 2975
rect 12069 2935 12127 2941
rect 12176 2944 12357 2972
rect 11330 2864 11336 2916
rect 11388 2904 11394 2916
rect 12176 2904 12204 2944
rect 12345 2941 12357 2944
rect 12391 2972 12403 2975
rect 16022 2972 16028 2984
rect 12391 2944 16028 2972
rect 12391 2941 12403 2944
rect 12345 2935 12403 2941
rect 16022 2932 16028 2944
rect 16080 2972 16086 2984
rect 17405 2975 17463 2981
rect 17405 2972 17417 2975
rect 16080 2944 17417 2972
rect 16080 2932 16086 2944
rect 17405 2941 17417 2944
rect 17451 2941 17463 2975
rect 17405 2935 17463 2941
rect 11388 2876 12204 2904
rect 11388 2864 11394 2876
rect 1486 2796 1492 2848
rect 1544 2796 1550 2848
rect 4430 2796 4436 2848
rect 4488 2836 4494 2848
rect 4985 2839 5043 2845
rect 4985 2836 4997 2839
rect 4488 2808 4997 2836
rect 4488 2796 4494 2808
rect 4985 2805 4997 2808
rect 5031 2805 5043 2839
rect 4985 2799 5043 2805
rect 8389 2839 8447 2845
rect 8389 2805 8401 2839
rect 8435 2836 8447 2839
rect 8662 2836 8668 2848
rect 8435 2808 8668 2836
rect 8435 2805 8447 2808
rect 8389 2799 8447 2805
rect 8662 2796 8668 2808
rect 8720 2796 8726 2848
rect 11103 2839 11161 2845
rect 11103 2805 11115 2839
rect 11149 2836 11161 2839
rect 11238 2836 11244 2848
rect 11149 2808 11244 2836
rect 11149 2805 11161 2808
rect 11103 2799 11161 2805
rect 11238 2796 11244 2808
rect 11296 2796 11302 2848
rect 18831 2839 18889 2845
rect 18831 2805 18843 2839
rect 18877 2836 18889 2839
rect 18966 2836 18972 2848
rect 18877 2808 18972 2836
rect 18877 2805 18889 2808
rect 18831 2799 18889 2805
rect 18966 2796 18972 2808
rect 19024 2796 19030 2848
rect 20162 2796 20168 2848
rect 20220 2796 20226 2848
rect 1104 2746 20700 2768
rect 1104 2694 3399 2746
rect 3451 2694 3463 2746
rect 3515 2694 3527 2746
rect 3579 2694 3591 2746
rect 3643 2694 3655 2746
rect 3707 2694 8298 2746
rect 8350 2694 8362 2746
rect 8414 2694 8426 2746
rect 8478 2694 8490 2746
rect 8542 2694 8554 2746
rect 8606 2694 13197 2746
rect 13249 2694 13261 2746
rect 13313 2694 13325 2746
rect 13377 2694 13389 2746
rect 13441 2694 13453 2746
rect 13505 2694 18096 2746
rect 18148 2694 18160 2746
rect 18212 2694 18224 2746
rect 18276 2694 18288 2746
rect 18340 2694 18352 2746
rect 18404 2694 20700 2746
rect 1104 2672 20700 2694
rect 10318 2592 10324 2644
rect 10376 2632 10382 2644
rect 10735 2635 10793 2641
rect 10735 2632 10747 2635
rect 10376 2604 10747 2632
rect 10376 2592 10382 2604
rect 10735 2601 10747 2604
rect 10781 2601 10793 2635
rect 10735 2595 10793 2601
rect 10594 2524 10600 2576
rect 10652 2564 10658 2576
rect 11057 2567 11115 2573
rect 11057 2564 11069 2567
rect 10652 2536 11069 2564
rect 10652 2524 10658 2536
rect 11057 2533 11069 2536
rect 11103 2533 11115 2567
rect 11057 2527 11115 2533
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 4982 2496 4988 2508
rect 4111 2468 4988 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 4982 2456 4988 2468
rect 5040 2456 5046 2508
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2465 5871 2499
rect 5813 2459 5871 2465
rect 1394 2388 1400 2440
rect 1452 2428 1458 2440
rect 1489 2431 1547 2437
rect 1489 2428 1501 2431
rect 1452 2400 1501 2428
rect 1452 2388 1458 2400
rect 1489 2397 1501 2400
rect 1535 2397 1547 2431
rect 1489 2391 1547 2397
rect 1946 2388 1952 2440
rect 2004 2388 2010 2440
rect 3234 2388 3240 2440
rect 3292 2388 3298 2440
rect 5828 2428 5856 2459
rect 8938 2456 8944 2508
rect 8996 2456 9002 2508
rect 9309 2499 9367 2505
rect 9309 2465 9321 2499
rect 9355 2496 9367 2499
rect 9490 2496 9496 2508
rect 9355 2468 9496 2496
rect 9355 2465 9367 2468
rect 9309 2459 9367 2465
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5828 2400 5917 2428
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 7098 2388 7104 2440
rect 7156 2388 7162 2440
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2428 8447 2431
rect 8662 2428 8668 2440
rect 8435 2400 8668 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 11238 2388 11244 2440
rect 11296 2388 11302 2440
rect 12526 2388 12532 2440
rect 12584 2388 12590 2440
rect 13538 2388 13544 2440
rect 13596 2388 13602 2440
rect 15010 2388 15016 2440
rect 15068 2428 15074 2440
rect 15105 2431 15163 2437
rect 15105 2428 15117 2431
rect 15068 2400 15117 2428
rect 15068 2388 15074 2400
rect 15105 2397 15117 2400
rect 15151 2397 15163 2431
rect 15105 2391 15163 2397
rect 16114 2388 16120 2440
rect 16172 2388 16178 2440
rect 17402 2388 17408 2440
rect 17460 2388 17466 2440
rect 18966 2388 18972 2440
rect 19024 2388 19030 2440
rect 19518 2388 19524 2440
rect 19576 2388 19582 2440
rect 20257 2431 20315 2437
rect 20257 2397 20269 2431
rect 20303 2428 20315 2431
rect 20438 2428 20444 2440
rect 20303 2400 20444 2428
rect 20303 2397 20315 2400
rect 20257 2391 20315 2397
rect 20438 2388 20444 2400
rect 20496 2388 20502 2440
rect 4341 2363 4399 2369
rect 4341 2329 4353 2363
rect 4387 2329 4399 2363
rect 4341 2323 4399 2329
rect 566 2252 572 2304
rect 624 2292 630 2304
rect 1581 2295 1639 2301
rect 1581 2292 1593 2295
rect 624 2264 1593 2292
rect 624 2252 630 2264
rect 1581 2261 1593 2264
rect 1627 2261 1639 2295
rect 1581 2255 1639 2261
rect 1854 2252 1860 2304
rect 1912 2292 1918 2304
rect 2133 2295 2191 2301
rect 2133 2292 2145 2295
rect 1912 2264 2145 2292
rect 1912 2252 1918 2264
rect 2133 2261 2145 2264
rect 2179 2261 2191 2295
rect 2133 2255 2191 2261
rect 3142 2252 3148 2304
rect 3200 2292 3206 2304
rect 3421 2295 3479 2301
rect 3421 2292 3433 2295
rect 3200 2264 3433 2292
rect 3200 2252 3206 2264
rect 3421 2261 3433 2264
rect 3467 2261 3479 2295
rect 4356 2292 4384 2323
rect 4798 2320 4804 2372
rect 4856 2320 4862 2372
rect 10502 2360 10508 2372
rect 10350 2332 10508 2360
rect 10502 2320 10508 2332
rect 10560 2320 10566 2372
rect 5258 2292 5264 2304
rect 4356 2264 5264 2292
rect 3421 2255 3479 2261
rect 5258 2252 5264 2264
rect 5316 2252 5322 2304
rect 5718 2252 5724 2304
rect 5776 2292 5782 2304
rect 6089 2295 6147 2301
rect 6089 2292 6101 2295
rect 5776 2264 6101 2292
rect 5776 2252 5782 2264
rect 6089 2261 6101 2264
rect 6135 2261 6147 2295
rect 6089 2255 6147 2261
rect 7006 2252 7012 2304
rect 7064 2292 7070 2304
rect 7285 2295 7343 2301
rect 7285 2292 7297 2295
rect 7064 2264 7297 2292
rect 7064 2252 7070 2264
rect 7285 2261 7297 2264
rect 7331 2261 7343 2295
rect 7285 2255 7343 2261
rect 8294 2252 8300 2304
rect 8352 2292 8358 2304
rect 8573 2295 8631 2301
rect 8573 2292 8585 2295
rect 8352 2264 8585 2292
rect 8352 2252 8358 2264
rect 8573 2261 8585 2264
rect 8619 2261 8631 2295
rect 8573 2255 8631 2261
rect 12158 2252 12164 2304
rect 12216 2292 12222 2304
rect 12345 2295 12403 2301
rect 12345 2292 12357 2295
rect 12216 2264 12357 2292
rect 12216 2252 12222 2264
rect 12345 2261 12357 2264
rect 12391 2261 12403 2295
rect 12345 2255 12403 2261
rect 13446 2252 13452 2304
rect 13504 2292 13510 2304
rect 13725 2295 13783 2301
rect 13725 2292 13737 2295
rect 13504 2264 13737 2292
rect 13504 2252 13510 2264
rect 13725 2261 13737 2264
rect 13771 2261 13783 2295
rect 13725 2255 13783 2261
rect 14734 2252 14740 2304
rect 14792 2292 14798 2304
rect 14921 2295 14979 2301
rect 14921 2292 14933 2295
rect 14792 2264 14933 2292
rect 14792 2252 14798 2264
rect 14921 2261 14933 2264
rect 14967 2261 14979 2295
rect 14921 2255 14979 2261
rect 16022 2252 16028 2304
rect 16080 2292 16086 2304
rect 16301 2295 16359 2301
rect 16301 2292 16313 2295
rect 16080 2264 16313 2292
rect 16080 2252 16086 2264
rect 16301 2261 16313 2264
rect 16347 2261 16359 2295
rect 16301 2255 16359 2261
rect 17310 2252 17316 2304
rect 17368 2292 17374 2304
rect 17589 2295 17647 2301
rect 17589 2292 17601 2295
rect 17368 2264 17601 2292
rect 17368 2252 17374 2264
rect 17589 2261 17601 2264
rect 17635 2261 17647 2295
rect 17589 2255 17647 2261
rect 18598 2252 18604 2304
rect 18656 2292 18662 2304
rect 18785 2295 18843 2301
rect 18785 2292 18797 2295
rect 18656 2264 18797 2292
rect 18656 2252 18662 2264
rect 18785 2261 18797 2264
rect 18831 2261 18843 2295
rect 18785 2255 18843 2261
rect 19705 2295 19763 2301
rect 19705 2261 19717 2295
rect 19751 2292 19763 2295
rect 19886 2292 19892 2304
rect 19751 2264 19892 2292
rect 19751 2261 19763 2264
rect 19705 2255 19763 2261
rect 19886 2252 19892 2264
rect 19944 2252 19950 2304
rect 20165 2295 20223 2301
rect 20165 2261 20177 2295
rect 20211 2292 20223 2295
rect 21174 2292 21180 2304
rect 20211 2264 21180 2292
rect 20211 2261 20223 2264
rect 20165 2255 20223 2261
rect 21174 2252 21180 2264
rect 21232 2252 21238 2304
rect 1104 2202 20859 2224
rect 1104 2150 5848 2202
rect 5900 2150 5912 2202
rect 5964 2150 5976 2202
rect 6028 2150 6040 2202
rect 6092 2150 6104 2202
rect 6156 2150 10747 2202
rect 10799 2150 10811 2202
rect 10863 2150 10875 2202
rect 10927 2150 10939 2202
rect 10991 2150 11003 2202
rect 11055 2150 15646 2202
rect 15698 2150 15710 2202
rect 15762 2150 15774 2202
rect 15826 2150 15838 2202
rect 15890 2150 15902 2202
rect 15954 2150 20545 2202
rect 20597 2150 20609 2202
rect 20661 2150 20673 2202
rect 20725 2150 20737 2202
rect 20789 2150 20801 2202
rect 20853 2150 20859 2202
rect 1104 2128 20859 2150
<< via1 >>
rect 5848 21734 5900 21786
rect 5912 21734 5964 21786
rect 5976 21734 6028 21786
rect 6040 21734 6092 21786
rect 6104 21734 6156 21786
rect 10747 21734 10799 21786
rect 10811 21734 10863 21786
rect 10875 21734 10927 21786
rect 10939 21734 10991 21786
rect 11003 21734 11055 21786
rect 15646 21734 15698 21786
rect 15710 21734 15762 21786
rect 15774 21734 15826 21786
rect 15838 21734 15890 21786
rect 15902 21734 15954 21786
rect 20545 21734 20597 21786
rect 20609 21734 20661 21786
rect 20673 21734 20725 21786
rect 20737 21734 20789 21786
rect 20801 21734 20853 21786
rect 572 21632 624 21684
rect 3148 21632 3200 21684
rect 5724 21632 5776 21684
rect 7012 21632 7064 21684
rect 8300 21632 8352 21684
rect 10600 21632 10652 21684
rect 13452 21632 13504 21684
rect 14740 21632 14792 21684
rect 16028 21632 16080 21684
rect 17592 21675 17644 21684
rect 17592 21641 17601 21675
rect 17601 21641 17635 21675
rect 17635 21641 17644 21675
rect 17592 21632 17644 21641
rect 18604 21632 18656 21684
rect 20076 21675 20128 21684
rect 20076 21641 20085 21675
rect 20085 21641 20119 21675
rect 20119 21641 20128 21675
rect 20076 21632 20128 21641
rect 1952 21607 2004 21616
rect 1952 21573 1961 21607
rect 1961 21573 1995 21607
rect 1995 21573 2004 21607
rect 1952 21564 2004 21573
rect 4528 21607 4580 21616
rect 4528 21573 4537 21607
rect 4537 21573 4571 21607
rect 4571 21573 4580 21607
rect 4528 21564 4580 21573
rect 9588 21564 9640 21616
rect 12164 21564 12216 21616
rect 1492 21539 1544 21548
rect 1492 21505 1501 21539
rect 1501 21505 1535 21539
rect 1535 21505 1544 21539
rect 1492 21496 1544 21505
rect 3056 21496 3108 21548
rect 3792 21496 3844 21548
rect 4896 21539 4948 21548
rect 4896 21505 4905 21539
rect 4905 21505 4939 21539
rect 4939 21505 4948 21539
rect 4896 21496 4948 21505
rect 5632 21496 5684 21548
rect 7196 21539 7248 21548
rect 7196 21505 7205 21539
rect 7205 21505 7239 21539
rect 7239 21505 7248 21539
rect 7196 21496 7248 21505
rect 8852 21496 8904 21548
rect 10048 21539 10100 21548
rect 10048 21505 10057 21539
rect 10057 21505 10091 21539
rect 10091 21505 10100 21539
rect 10048 21496 10100 21505
rect 11612 21539 11664 21548
rect 11612 21505 11621 21539
rect 11621 21505 11655 21539
rect 11655 21505 11664 21539
rect 11612 21496 11664 21505
rect 12624 21539 12676 21548
rect 12624 21505 12633 21539
rect 12633 21505 12667 21539
rect 12667 21505 12676 21539
rect 12624 21496 12676 21505
rect 14188 21539 14240 21548
rect 14188 21505 14197 21539
rect 14197 21505 14231 21539
rect 14231 21505 14240 21539
rect 14188 21496 14240 21505
rect 15016 21496 15068 21548
rect 16764 21539 16816 21548
rect 16764 21505 16773 21539
rect 16773 21505 16807 21539
rect 16807 21505 16816 21539
rect 16764 21496 16816 21505
rect 17500 21539 17552 21548
rect 17500 21505 17509 21539
rect 17509 21505 17543 21539
rect 17543 21505 17552 21539
rect 17500 21496 17552 21505
rect 19340 21539 19392 21548
rect 19340 21505 19349 21539
rect 19349 21505 19383 21539
rect 19383 21505 19392 21539
rect 19340 21496 19392 21505
rect 19708 21496 19760 21548
rect 3399 21190 3451 21242
rect 3463 21190 3515 21242
rect 3527 21190 3579 21242
rect 3591 21190 3643 21242
rect 3655 21190 3707 21242
rect 8298 21190 8350 21242
rect 8362 21190 8414 21242
rect 8426 21190 8478 21242
rect 8490 21190 8542 21242
rect 8554 21190 8606 21242
rect 13197 21190 13249 21242
rect 13261 21190 13313 21242
rect 13325 21190 13377 21242
rect 13389 21190 13441 21242
rect 13453 21190 13505 21242
rect 18096 21190 18148 21242
rect 18160 21190 18212 21242
rect 18224 21190 18276 21242
rect 18288 21190 18340 21242
rect 18352 21190 18404 21242
rect 1308 21088 1360 21140
rect 8944 20952 8996 21004
rect 3976 20859 4028 20868
rect 3976 20825 3985 20859
rect 3985 20825 4019 20859
rect 4019 20825 4028 20859
rect 3976 20816 4028 20825
rect 4804 20927 4856 20936
rect 4804 20893 4813 20927
rect 4813 20893 4847 20927
rect 4847 20893 4856 20927
rect 4804 20884 4856 20893
rect 7288 20927 7340 20936
rect 7288 20893 7297 20927
rect 7297 20893 7331 20927
rect 7331 20893 7340 20927
rect 7288 20884 7340 20893
rect 8208 20884 8260 20936
rect 9772 20884 9824 20936
rect 12624 21088 12676 21140
rect 19340 21088 19392 21140
rect 21180 21088 21232 21140
rect 15384 20952 15436 21004
rect 6736 20816 6788 20868
rect 7840 20859 7892 20868
rect 7840 20825 7849 20859
rect 7849 20825 7883 20859
rect 7883 20825 7892 20859
rect 7840 20816 7892 20825
rect 9312 20859 9364 20868
rect 9312 20825 9321 20859
rect 9321 20825 9355 20859
rect 9355 20825 9364 20859
rect 9312 20816 9364 20825
rect 5080 20748 5132 20800
rect 9036 20791 9088 20800
rect 9036 20757 9045 20791
rect 9045 20757 9079 20791
rect 9079 20757 9088 20791
rect 9036 20748 9088 20757
rect 9588 20748 9640 20800
rect 10508 20748 10560 20800
rect 12532 20816 12584 20868
rect 13084 20816 13136 20868
rect 17040 20927 17092 20936
rect 17040 20893 17049 20927
rect 17049 20893 17083 20927
rect 17083 20893 17092 20927
rect 17040 20884 17092 20893
rect 19616 20927 19668 20936
rect 19616 20893 19625 20927
rect 19625 20893 19659 20927
rect 19659 20893 19668 20927
rect 19616 20884 19668 20893
rect 13820 20859 13872 20868
rect 13820 20825 13829 20859
rect 13829 20825 13863 20859
rect 13863 20825 13872 20859
rect 13820 20816 13872 20825
rect 14372 20859 14424 20868
rect 14372 20825 14381 20859
rect 14381 20825 14415 20859
rect 14415 20825 14424 20859
rect 14372 20816 14424 20825
rect 15200 20748 15252 20800
rect 18972 20816 19024 20868
rect 20168 20816 20220 20868
rect 20260 20859 20312 20868
rect 20260 20825 20269 20859
rect 20269 20825 20303 20859
rect 20303 20825 20312 20859
rect 20260 20816 20312 20825
rect 19432 20748 19484 20800
rect 5848 20646 5900 20698
rect 5912 20646 5964 20698
rect 5976 20646 6028 20698
rect 6040 20646 6092 20698
rect 6104 20646 6156 20698
rect 10747 20646 10799 20698
rect 10811 20646 10863 20698
rect 10875 20646 10927 20698
rect 10939 20646 10991 20698
rect 11003 20646 11055 20698
rect 15646 20646 15698 20698
rect 15710 20646 15762 20698
rect 15774 20646 15826 20698
rect 15838 20646 15890 20698
rect 15902 20646 15954 20698
rect 20545 20646 20597 20698
rect 20609 20646 20661 20698
rect 20673 20646 20725 20698
rect 20737 20646 20789 20698
rect 20801 20646 20853 20698
rect 11612 20544 11664 20596
rect 14372 20544 14424 20596
rect 20260 20544 20312 20596
rect 6736 20476 6788 20528
rect 9036 20476 9088 20528
rect 9956 20476 10008 20528
rect 12808 20476 12860 20528
rect 19616 20476 19668 20528
rect 9588 20451 9640 20460
rect 9588 20417 9597 20451
rect 9597 20417 9631 20451
rect 9631 20417 9640 20451
rect 9588 20408 9640 20417
rect 18328 20451 18380 20460
rect 18328 20417 18372 20451
rect 18372 20417 18380 20451
rect 18328 20408 18380 20417
rect 4252 20340 4304 20392
rect 5080 20340 5132 20392
rect 7012 20340 7064 20392
rect 7288 20340 7340 20392
rect 7656 20383 7708 20392
rect 7656 20349 7665 20383
rect 7665 20349 7699 20383
rect 7699 20349 7708 20383
rect 7656 20340 7708 20349
rect 9404 20340 9456 20392
rect 11520 20340 11572 20392
rect 13084 20383 13136 20392
rect 13084 20349 13093 20383
rect 13093 20349 13127 20383
rect 13127 20349 13136 20383
rect 13084 20340 13136 20349
rect 13912 20340 13964 20392
rect 17960 20340 18012 20392
rect 4068 20204 4120 20256
rect 5356 20247 5408 20256
rect 5356 20213 5365 20247
rect 5365 20213 5399 20247
rect 5399 20213 5408 20247
rect 5356 20204 5408 20213
rect 9128 20247 9180 20256
rect 9128 20213 9137 20247
rect 9137 20213 9171 20247
rect 9171 20213 9180 20247
rect 9128 20204 9180 20213
rect 16488 20204 16540 20256
rect 16672 20204 16724 20256
rect 3399 20102 3451 20154
rect 3463 20102 3515 20154
rect 3527 20102 3579 20154
rect 3591 20102 3643 20154
rect 3655 20102 3707 20154
rect 8298 20102 8350 20154
rect 8362 20102 8414 20154
rect 8426 20102 8478 20154
rect 8490 20102 8542 20154
rect 8554 20102 8606 20154
rect 13197 20102 13249 20154
rect 13261 20102 13313 20154
rect 13325 20102 13377 20154
rect 13389 20102 13441 20154
rect 13453 20102 13505 20154
rect 18096 20102 18148 20154
rect 18160 20102 18212 20154
rect 18224 20102 18276 20154
rect 18288 20102 18340 20154
rect 18352 20102 18404 20154
rect 4804 20000 4856 20052
rect 7656 20000 7708 20052
rect 8944 20000 8996 20052
rect 13912 20043 13964 20052
rect 13912 20009 13921 20043
rect 13921 20009 13955 20043
rect 13955 20009 13964 20043
rect 13912 20000 13964 20009
rect 17500 20000 17552 20052
rect 15200 19864 15252 19916
rect 4252 19796 4304 19848
rect 8392 19839 8444 19848
rect 8392 19805 8401 19839
rect 8401 19805 8435 19839
rect 8435 19805 8444 19839
rect 8392 19796 8444 19805
rect 9128 19839 9180 19848
rect 9128 19805 9136 19839
rect 9136 19805 9180 19839
rect 9128 19796 9180 19805
rect 11520 19796 11572 19848
rect 15292 19839 15344 19848
rect 15292 19805 15336 19839
rect 15336 19805 15344 19839
rect 15292 19796 15344 19805
rect 8944 19728 8996 19780
rect 12440 19771 12492 19780
rect 12440 19737 12449 19771
rect 12449 19737 12483 19771
rect 12483 19737 12492 19771
rect 12440 19728 12492 19737
rect 15568 19839 15620 19848
rect 15568 19805 15577 19839
rect 15577 19805 15611 19839
rect 15611 19805 15620 19839
rect 15568 19796 15620 19805
rect 18420 19796 18472 19848
rect 20352 19839 20404 19848
rect 20352 19805 20361 19839
rect 20361 19805 20395 19839
rect 20395 19805 20404 19839
rect 20352 19796 20404 19805
rect 16672 19728 16724 19780
rect 12808 19660 12860 19712
rect 13820 19660 13872 19712
rect 18236 19660 18288 19712
rect 5848 19558 5900 19610
rect 5912 19558 5964 19610
rect 5976 19558 6028 19610
rect 6040 19558 6092 19610
rect 6104 19558 6156 19610
rect 10747 19558 10799 19610
rect 10811 19558 10863 19610
rect 10875 19558 10927 19610
rect 10939 19558 10991 19610
rect 11003 19558 11055 19610
rect 15646 19558 15698 19610
rect 15710 19558 15762 19610
rect 15774 19558 15826 19610
rect 15838 19558 15890 19610
rect 15902 19558 15954 19610
rect 20545 19558 20597 19610
rect 20609 19558 20661 19610
rect 20673 19558 20725 19610
rect 20737 19558 20789 19610
rect 20801 19558 20853 19610
rect 1492 19456 1544 19508
rect 4344 19456 4396 19508
rect 2136 19388 2188 19440
rect 2964 19388 3016 19440
rect 6736 19456 6788 19508
rect 12440 19456 12492 19508
rect 19708 19499 19760 19508
rect 19708 19465 19717 19499
rect 19717 19465 19751 19499
rect 19751 19465 19760 19499
rect 19708 19456 19760 19465
rect 5356 19388 5408 19440
rect 9036 19388 9088 19440
rect 12808 19388 12860 19440
rect 18236 19431 18288 19440
rect 18236 19397 18245 19431
rect 18245 19397 18279 19431
rect 18279 19397 18288 19431
rect 18236 19388 18288 19397
rect 18788 19388 18840 19440
rect 7840 19320 7892 19372
rect 8024 19320 8076 19372
rect 10324 19320 10376 19372
rect 11520 19363 11572 19372
rect 11520 19329 11529 19363
rect 11529 19329 11563 19363
rect 11563 19329 11572 19363
rect 11520 19320 11572 19329
rect 17960 19363 18012 19372
rect 17960 19329 17969 19363
rect 17969 19329 18003 19363
rect 18003 19329 18012 19363
rect 17960 19320 18012 19329
rect 2872 19295 2924 19304
rect 2872 19261 2881 19295
rect 2881 19261 2915 19295
rect 2915 19261 2924 19295
rect 2872 19252 2924 19261
rect 8852 19252 8904 19304
rect 11796 19295 11848 19304
rect 11796 19261 11805 19295
rect 11805 19261 11839 19295
rect 11839 19261 11848 19295
rect 11796 19252 11848 19261
rect 5172 19116 5224 19168
rect 9680 19116 9732 19168
rect 3399 19014 3451 19066
rect 3463 19014 3515 19066
rect 3527 19014 3579 19066
rect 3591 19014 3643 19066
rect 3655 19014 3707 19066
rect 8298 19014 8350 19066
rect 8362 19014 8414 19066
rect 8426 19014 8478 19066
rect 8490 19014 8542 19066
rect 8554 19014 8606 19066
rect 13197 19014 13249 19066
rect 13261 19014 13313 19066
rect 13325 19014 13377 19066
rect 13389 19014 13441 19066
rect 13453 19014 13505 19066
rect 18096 19014 18148 19066
rect 18160 19014 18212 19066
rect 18224 19014 18276 19066
rect 18288 19014 18340 19066
rect 18352 19014 18404 19066
rect 2872 18912 2924 18964
rect 11796 18912 11848 18964
rect 8024 18776 8076 18828
rect 10324 18819 10376 18828
rect 10324 18785 10333 18819
rect 10333 18785 10367 18819
rect 10367 18785 10376 18819
rect 10324 18776 10376 18785
rect 1952 18751 2004 18760
rect 1952 18717 1970 18751
rect 1970 18717 2004 18751
rect 1952 18708 2004 18717
rect 4068 18708 4120 18760
rect 5172 18751 5224 18760
rect 5172 18717 5181 18751
rect 5181 18717 5215 18751
rect 5215 18717 5224 18751
rect 5172 18708 5224 18717
rect 16028 18708 16080 18760
rect 17592 18751 17644 18760
rect 17592 18717 17601 18751
rect 17601 18717 17635 18751
rect 17635 18717 17644 18751
rect 17592 18708 17644 18717
rect 18788 18708 18840 18760
rect 20076 18751 20128 18760
rect 20076 18717 20085 18751
rect 20085 18717 20119 18751
rect 20119 18717 20128 18751
rect 20076 18708 20128 18717
rect 5724 18640 5776 18692
rect 6736 18640 6788 18692
rect 10600 18683 10652 18692
rect 10600 18649 10609 18683
rect 10609 18649 10643 18683
rect 10643 18649 10652 18683
rect 10600 18640 10652 18649
rect 6920 18615 6972 18624
rect 6920 18581 6929 18615
rect 6929 18581 6963 18615
rect 6963 18581 6972 18615
rect 6920 18572 6972 18581
rect 9312 18572 9364 18624
rect 12808 18572 12860 18624
rect 20260 18615 20312 18624
rect 20260 18581 20269 18615
rect 20269 18581 20303 18615
rect 20303 18581 20312 18615
rect 20260 18572 20312 18581
rect 5848 18470 5900 18522
rect 5912 18470 5964 18522
rect 5976 18470 6028 18522
rect 6040 18470 6092 18522
rect 6104 18470 6156 18522
rect 10747 18470 10799 18522
rect 10811 18470 10863 18522
rect 10875 18470 10927 18522
rect 10939 18470 10991 18522
rect 11003 18470 11055 18522
rect 15646 18470 15698 18522
rect 15710 18470 15762 18522
rect 15774 18470 15826 18522
rect 15838 18470 15890 18522
rect 15902 18470 15954 18522
rect 20545 18470 20597 18522
rect 20609 18470 20661 18522
rect 20673 18470 20725 18522
rect 20737 18470 20789 18522
rect 20801 18470 20853 18522
rect 5724 18368 5776 18420
rect 8852 18368 8904 18420
rect 9312 18368 9364 18420
rect 4344 18343 4396 18352
rect 4344 18309 4353 18343
rect 4353 18309 4387 18343
rect 4387 18309 4396 18343
rect 4344 18300 4396 18309
rect 6736 18300 6788 18352
rect 9036 18300 9088 18352
rect 9680 18300 9732 18352
rect 10600 18368 10652 18420
rect 16028 18411 16080 18420
rect 16028 18377 16037 18411
rect 16037 18377 16071 18411
rect 16071 18377 16080 18411
rect 16028 18368 16080 18377
rect 14372 18275 14424 18284
rect 14372 18241 14381 18275
rect 14381 18241 14415 18275
rect 14415 18241 14424 18275
rect 14372 18232 14424 18241
rect 15660 18300 15712 18352
rect 18420 18300 18472 18352
rect 18788 18300 18840 18352
rect 4068 18207 4120 18216
rect 4068 18173 4077 18207
rect 4077 18173 4111 18207
rect 4111 18173 4120 18207
rect 4068 18164 4120 18173
rect 7012 18207 7064 18216
rect 7012 18173 7021 18207
rect 7021 18173 7055 18207
rect 7055 18173 7064 18207
rect 7012 18164 7064 18173
rect 7840 18164 7892 18216
rect 8024 18164 8076 18216
rect 17868 18275 17920 18284
rect 17868 18241 17877 18275
rect 17877 18241 17911 18275
rect 17911 18241 17920 18275
rect 17868 18232 17920 18241
rect 15660 18139 15712 18148
rect 15660 18105 15669 18139
rect 15669 18105 15703 18139
rect 15703 18105 15712 18139
rect 15660 18096 15712 18105
rect 15292 18028 15344 18080
rect 15568 18071 15620 18080
rect 15568 18037 15577 18071
rect 15577 18037 15611 18071
rect 15611 18037 15620 18071
rect 15568 18028 15620 18037
rect 19524 18028 19576 18080
rect 3399 17926 3451 17978
rect 3463 17926 3515 17978
rect 3527 17926 3579 17978
rect 3591 17926 3643 17978
rect 3655 17926 3707 17978
rect 8298 17926 8350 17978
rect 8362 17926 8414 17978
rect 8426 17926 8478 17978
rect 8490 17926 8542 17978
rect 8554 17926 8606 17978
rect 13197 17926 13249 17978
rect 13261 17926 13313 17978
rect 13325 17926 13377 17978
rect 13389 17926 13441 17978
rect 13453 17926 13505 17978
rect 18096 17926 18148 17978
rect 18160 17926 18212 17978
rect 18224 17926 18276 17978
rect 18288 17926 18340 17978
rect 18352 17926 18404 17978
rect 3792 17824 3844 17876
rect 1492 17663 1544 17672
rect 1492 17629 1501 17663
rect 1501 17629 1535 17663
rect 1535 17629 1544 17663
rect 1492 17620 1544 17629
rect 1860 17663 1912 17672
rect 1860 17629 1869 17663
rect 1869 17629 1903 17663
rect 1903 17629 1912 17663
rect 1860 17620 1912 17629
rect 4068 17620 4120 17672
rect 7012 17824 7064 17876
rect 7840 17867 7892 17876
rect 7840 17833 7849 17867
rect 7849 17833 7883 17867
rect 7883 17833 7892 17867
rect 7840 17824 7892 17833
rect 9956 17824 10008 17876
rect 6920 17688 6972 17740
rect 13728 17688 13780 17740
rect 13544 17663 13596 17672
rect 2872 17552 2924 17604
rect 2136 17484 2188 17536
rect 3516 17484 3568 17536
rect 6736 17484 6788 17536
rect 9036 17552 9088 17604
rect 13544 17629 13553 17663
rect 13553 17629 13587 17663
rect 13587 17629 13596 17663
rect 13544 17620 13596 17629
rect 14096 17663 14148 17672
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 15660 17824 15712 17876
rect 19616 17867 19668 17876
rect 19616 17833 19625 17867
rect 19625 17833 19659 17867
rect 19659 17833 19668 17867
rect 19616 17824 19668 17833
rect 20076 17824 20128 17876
rect 17592 17688 17644 17740
rect 16488 17620 16540 17672
rect 18052 17620 18104 17672
rect 12532 17552 12584 17604
rect 18512 17552 18564 17604
rect 20076 17663 20128 17672
rect 20076 17629 20085 17663
rect 20085 17629 20119 17663
rect 20119 17629 20128 17663
rect 20076 17620 20128 17629
rect 11244 17484 11296 17536
rect 17960 17484 18012 17536
rect 20260 17527 20312 17536
rect 20260 17493 20269 17527
rect 20269 17493 20303 17527
rect 20303 17493 20312 17527
rect 20260 17484 20312 17493
rect 5848 17382 5900 17434
rect 5912 17382 5964 17434
rect 5976 17382 6028 17434
rect 6040 17382 6092 17434
rect 6104 17382 6156 17434
rect 10747 17382 10799 17434
rect 10811 17382 10863 17434
rect 10875 17382 10927 17434
rect 10939 17382 10991 17434
rect 11003 17382 11055 17434
rect 15646 17382 15698 17434
rect 15710 17382 15762 17434
rect 15774 17382 15826 17434
rect 15838 17382 15890 17434
rect 15902 17382 15954 17434
rect 20545 17382 20597 17434
rect 20609 17382 20661 17434
rect 20673 17382 20725 17434
rect 20737 17382 20789 17434
rect 20801 17382 20853 17434
rect 1860 17280 1912 17332
rect 2872 17280 2924 17332
rect 10048 17280 10100 17332
rect 11244 17280 11296 17332
rect 14372 17280 14424 17332
rect 17040 17280 17092 17332
rect 17224 17323 17276 17332
rect 17224 17289 17233 17323
rect 17233 17289 17267 17323
rect 17267 17289 17276 17323
rect 17224 17280 17276 17289
rect 18052 17323 18104 17332
rect 18052 17289 18061 17323
rect 18061 17289 18095 17323
rect 18095 17289 18104 17323
rect 18052 17280 18104 17289
rect 9956 17212 10008 17264
rect 13544 17212 13596 17264
rect 1952 17144 2004 17196
rect 3516 17187 3568 17196
rect 3516 17153 3525 17187
rect 3525 17153 3559 17187
rect 3559 17153 3568 17187
rect 3516 17144 3568 17153
rect 3792 17076 3844 17128
rect 9588 17144 9640 17196
rect 3148 16940 3200 16992
rect 3240 16940 3292 16992
rect 3976 16940 4028 16992
rect 9496 17076 9548 17128
rect 9772 17076 9824 17128
rect 14096 17144 14148 17196
rect 14924 17144 14976 17196
rect 17684 17212 17736 17264
rect 19616 17212 19668 17264
rect 15476 17144 15528 17196
rect 13728 17076 13780 17128
rect 9772 16940 9824 16992
rect 15660 16983 15712 16992
rect 15660 16949 15669 16983
rect 15669 16949 15703 16983
rect 15703 16949 15712 16983
rect 15660 16940 15712 16949
rect 17500 17187 17552 17196
rect 17500 17153 17509 17187
rect 17509 17153 17543 17187
rect 17543 17153 17552 17187
rect 17500 17144 17552 17153
rect 17960 17144 18012 17196
rect 17132 17008 17184 17060
rect 18420 16940 18472 16992
rect 20444 16940 20496 16992
rect 3399 16838 3451 16890
rect 3463 16838 3515 16890
rect 3527 16838 3579 16890
rect 3591 16838 3643 16890
rect 3655 16838 3707 16890
rect 8298 16838 8350 16890
rect 8362 16838 8414 16890
rect 8426 16838 8478 16890
rect 8490 16838 8542 16890
rect 8554 16838 8606 16890
rect 13197 16838 13249 16890
rect 13261 16838 13313 16890
rect 13325 16838 13377 16890
rect 13389 16838 13441 16890
rect 13453 16838 13505 16890
rect 18096 16838 18148 16890
rect 18160 16838 18212 16890
rect 18224 16838 18276 16890
rect 18288 16838 18340 16890
rect 18352 16838 18404 16890
rect 9588 16736 9640 16788
rect 12808 16736 12860 16788
rect 17132 16779 17184 16788
rect 17132 16745 17141 16779
rect 17141 16745 17175 16779
rect 17175 16745 17184 16779
rect 17132 16736 17184 16745
rect 17500 16736 17552 16788
rect 19892 16668 19944 16720
rect 2872 16600 2924 16652
rect 3240 16600 3292 16652
rect 3148 16575 3200 16584
rect 3148 16541 3157 16575
rect 3157 16541 3191 16575
rect 3191 16541 3200 16575
rect 3148 16532 3200 16541
rect 3792 16532 3844 16584
rect 9312 16600 9364 16652
rect 15384 16643 15436 16652
rect 15384 16609 15393 16643
rect 15393 16609 15427 16643
rect 15427 16609 15436 16643
rect 15384 16600 15436 16609
rect 15660 16643 15712 16652
rect 15660 16609 15669 16643
rect 15669 16609 15703 16643
rect 15703 16609 15712 16643
rect 15660 16600 15712 16609
rect 8024 16575 8076 16584
rect 8024 16541 8033 16575
rect 8033 16541 8067 16575
rect 8067 16541 8076 16575
rect 8024 16532 8076 16541
rect 9864 16532 9916 16584
rect 4988 16439 5040 16448
rect 4988 16405 4997 16439
rect 4997 16405 5031 16439
rect 5031 16405 5040 16439
rect 4988 16396 5040 16405
rect 16580 16396 16632 16448
rect 17132 16532 17184 16584
rect 19984 16464 20036 16516
rect 20168 16464 20220 16516
rect 17408 16396 17460 16448
rect 5848 16294 5900 16346
rect 5912 16294 5964 16346
rect 5976 16294 6028 16346
rect 6040 16294 6092 16346
rect 6104 16294 6156 16346
rect 10747 16294 10799 16346
rect 10811 16294 10863 16346
rect 10875 16294 10927 16346
rect 10939 16294 10991 16346
rect 11003 16294 11055 16346
rect 15646 16294 15698 16346
rect 15710 16294 15762 16346
rect 15774 16294 15826 16346
rect 15838 16294 15890 16346
rect 15902 16294 15954 16346
rect 20545 16294 20597 16346
rect 20609 16294 20661 16346
rect 20673 16294 20725 16346
rect 20737 16294 20789 16346
rect 20801 16294 20853 16346
rect 9864 16235 9916 16244
rect 9864 16201 9873 16235
rect 9873 16201 9907 16235
rect 9907 16201 9916 16235
rect 9864 16192 9916 16201
rect 20076 16192 20128 16244
rect 7840 16124 7892 16176
rect 17960 16124 18012 16176
rect 6184 16056 6236 16108
rect 8024 15988 8076 16040
rect 9220 15988 9272 16040
rect 11244 16056 11296 16108
rect 19892 16056 19944 16108
rect 18512 16031 18564 16040
rect 18512 15997 18521 16031
rect 18521 15997 18555 16031
rect 18555 15997 18564 16031
rect 18512 15988 18564 15997
rect 6368 15852 6420 15904
rect 14924 15852 14976 15904
rect 3399 15750 3451 15802
rect 3463 15750 3515 15802
rect 3527 15750 3579 15802
rect 3591 15750 3643 15802
rect 3655 15750 3707 15802
rect 8298 15750 8350 15802
rect 8362 15750 8414 15802
rect 8426 15750 8478 15802
rect 8490 15750 8542 15802
rect 8554 15750 8606 15802
rect 13197 15750 13249 15802
rect 13261 15750 13313 15802
rect 13325 15750 13377 15802
rect 13389 15750 13441 15802
rect 13453 15750 13505 15802
rect 18096 15750 18148 15802
rect 18160 15750 18212 15802
rect 18224 15750 18276 15802
rect 18288 15750 18340 15802
rect 18352 15750 18404 15802
rect 3056 15648 3108 15700
rect 3332 15648 3384 15700
rect 3976 15648 4028 15700
rect 11244 15691 11296 15700
rect 11244 15657 11253 15691
rect 11253 15657 11287 15691
rect 11287 15657 11296 15691
rect 11244 15648 11296 15657
rect 14188 15648 14240 15700
rect 15384 15648 15436 15700
rect 3240 15512 3292 15564
rect 9220 15555 9272 15564
rect 9220 15521 9229 15555
rect 9229 15521 9263 15555
rect 9263 15521 9272 15555
rect 9220 15512 9272 15521
rect 1768 15487 1820 15496
rect 1768 15453 1777 15487
rect 1777 15453 1811 15487
rect 1811 15453 1820 15487
rect 1768 15444 1820 15453
rect 3976 15487 4028 15496
rect 3976 15453 3984 15487
rect 3984 15453 4028 15487
rect 2688 15376 2740 15428
rect 3976 15444 4028 15453
rect 4988 15444 5040 15496
rect 7748 15444 7800 15496
rect 8392 15487 8444 15496
rect 8392 15453 8401 15487
rect 8401 15453 8435 15487
rect 8435 15453 8444 15487
rect 8392 15444 8444 15453
rect 3516 15308 3568 15360
rect 3976 15308 4028 15360
rect 7748 15308 7800 15360
rect 9680 15376 9732 15428
rect 8668 15308 8720 15360
rect 9956 15308 10008 15360
rect 11612 15487 11664 15496
rect 11612 15453 11621 15487
rect 11621 15453 11655 15487
rect 11655 15453 11664 15487
rect 11612 15444 11664 15453
rect 14372 15580 14424 15632
rect 14924 15555 14976 15564
rect 14924 15521 14933 15555
rect 14933 15521 14967 15555
rect 14967 15521 14976 15555
rect 14924 15512 14976 15521
rect 19340 15648 19392 15700
rect 19984 15648 20036 15700
rect 17132 15512 17184 15564
rect 12440 15376 12492 15428
rect 13268 15376 13320 15428
rect 14556 15376 14608 15428
rect 19800 15487 19852 15496
rect 19800 15453 19809 15487
rect 19809 15453 19843 15487
rect 19843 15453 19852 15487
rect 19800 15444 19852 15453
rect 14280 15308 14332 15360
rect 17500 15376 17552 15428
rect 19432 15376 19484 15428
rect 18512 15351 18564 15360
rect 18512 15317 18521 15351
rect 18521 15317 18555 15351
rect 18555 15317 18564 15351
rect 18512 15308 18564 15317
rect 19248 15308 19300 15360
rect 5848 15206 5900 15258
rect 5912 15206 5964 15258
rect 5976 15206 6028 15258
rect 6040 15206 6092 15258
rect 6104 15206 6156 15258
rect 10747 15206 10799 15258
rect 10811 15206 10863 15258
rect 10875 15206 10927 15258
rect 10939 15206 10991 15258
rect 11003 15206 11055 15258
rect 15646 15206 15698 15258
rect 15710 15206 15762 15258
rect 15774 15206 15826 15258
rect 15838 15206 15890 15258
rect 15902 15206 15954 15258
rect 20545 15206 20597 15258
rect 20609 15206 20661 15258
rect 20673 15206 20725 15258
rect 20737 15206 20789 15258
rect 20801 15206 20853 15258
rect 1768 15104 1820 15156
rect 2136 15104 2188 15156
rect 2688 15104 2740 15156
rect 4896 15104 4948 15156
rect 6184 15104 6236 15156
rect 7380 15104 7432 15156
rect 3332 14968 3384 15020
rect 3516 14968 3568 15020
rect 6368 15011 6420 15020
rect 6368 14977 6377 15011
rect 6377 14977 6411 15011
rect 6411 14977 6420 15011
rect 6368 14968 6420 14977
rect 7748 14968 7800 15020
rect 8024 15104 8076 15156
rect 8392 15147 8444 15156
rect 8392 15113 8401 15147
rect 8401 15113 8435 15147
rect 8435 15113 8444 15147
rect 8392 15104 8444 15113
rect 9772 15104 9824 15156
rect 9956 15036 10008 15088
rect 15016 15104 15068 15156
rect 17960 15104 18012 15156
rect 13268 15079 13320 15088
rect 13268 15045 13277 15079
rect 13277 15045 13311 15079
rect 13311 15045 13320 15079
rect 13268 15036 13320 15045
rect 14004 15036 14056 15088
rect 19800 15104 19852 15156
rect 19892 15036 19944 15088
rect 11152 14968 11204 15020
rect 18512 14968 18564 15020
rect 3056 14943 3108 14952
rect 3056 14909 3065 14943
rect 3065 14909 3099 14943
rect 3099 14909 3108 14943
rect 3056 14900 3108 14909
rect 5172 14900 5224 14952
rect 11612 14900 11664 14952
rect 13912 14900 13964 14952
rect 17684 14900 17736 14952
rect 18604 14943 18656 14952
rect 18604 14909 18613 14943
rect 18613 14909 18647 14943
rect 18647 14909 18656 14943
rect 18604 14900 18656 14909
rect 17040 14832 17092 14884
rect 11152 14807 11204 14816
rect 11152 14773 11161 14807
rect 11161 14773 11195 14807
rect 11195 14773 11204 14807
rect 11152 14764 11204 14773
rect 3399 14662 3451 14714
rect 3463 14662 3515 14714
rect 3527 14662 3579 14714
rect 3591 14662 3643 14714
rect 3655 14662 3707 14714
rect 8298 14662 8350 14714
rect 8362 14662 8414 14714
rect 8426 14662 8478 14714
rect 8490 14662 8542 14714
rect 8554 14662 8606 14714
rect 13197 14662 13249 14714
rect 13261 14662 13313 14714
rect 13325 14662 13377 14714
rect 13389 14662 13441 14714
rect 13453 14662 13505 14714
rect 18096 14662 18148 14714
rect 18160 14662 18212 14714
rect 18224 14662 18276 14714
rect 18288 14662 18340 14714
rect 18352 14662 18404 14714
rect 5172 14603 5224 14612
rect 5172 14569 5181 14603
rect 5181 14569 5215 14603
rect 5215 14569 5224 14603
rect 5172 14560 5224 14569
rect 16580 14560 16632 14612
rect 17040 14603 17092 14612
rect 17040 14569 17049 14603
rect 17049 14569 17083 14603
rect 17083 14569 17092 14603
rect 17040 14560 17092 14569
rect 17224 14492 17276 14544
rect 13912 14424 13964 14476
rect 17684 14424 17736 14476
rect 4988 14399 5040 14408
rect 4988 14365 4997 14399
rect 4997 14365 5031 14399
rect 5031 14365 5040 14399
rect 4988 14356 5040 14365
rect 17132 14356 17184 14408
rect 14280 14288 14332 14340
rect 15384 14288 15436 14340
rect 18420 14263 18472 14272
rect 18420 14229 18429 14263
rect 18429 14229 18463 14263
rect 18463 14229 18472 14263
rect 18420 14220 18472 14229
rect 5848 14118 5900 14170
rect 5912 14118 5964 14170
rect 5976 14118 6028 14170
rect 6040 14118 6092 14170
rect 6104 14118 6156 14170
rect 10747 14118 10799 14170
rect 10811 14118 10863 14170
rect 10875 14118 10927 14170
rect 10939 14118 10991 14170
rect 11003 14118 11055 14170
rect 15646 14118 15698 14170
rect 15710 14118 15762 14170
rect 15774 14118 15826 14170
rect 15838 14118 15890 14170
rect 15902 14118 15954 14170
rect 20545 14118 20597 14170
rect 20609 14118 20661 14170
rect 20673 14118 20725 14170
rect 20737 14118 20789 14170
rect 20801 14118 20853 14170
rect 8668 13948 8720 14000
rect 18420 13948 18472 14000
rect 19892 13948 19944 14000
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 2228 13923 2280 13932
rect 2228 13889 2237 13923
rect 2237 13889 2271 13923
rect 2271 13889 2280 13923
rect 2228 13880 2280 13889
rect 13084 13880 13136 13932
rect 3976 13855 4028 13864
rect 3976 13821 3985 13855
rect 3985 13821 4019 13855
rect 4019 13821 4028 13855
rect 3976 13812 4028 13821
rect 7840 13855 7892 13864
rect 7840 13821 7849 13855
rect 7849 13821 7883 13855
rect 7883 13821 7892 13855
rect 7840 13812 7892 13821
rect 1492 13676 1544 13728
rect 11152 13744 11204 13796
rect 12532 13744 12584 13796
rect 14556 13880 14608 13932
rect 15384 13812 15436 13864
rect 18604 13855 18656 13864
rect 18604 13821 18613 13855
rect 18613 13821 18647 13855
rect 18647 13821 18656 13855
rect 18604 13812 18656 13821
rect 9588 13719 9640 13728
rect 9588 13685 9597 13719
rect 9597 13685 9631 13719
rect 9631 13685 9640 13719
rect 9588 13676 9640 13685
rect 20352 13719 20404 13728
rect 20352 13685 20361 13719
rect 20361 13685 20395 13719
rect 20395 13685 20404 13719
rect 20352 13676 20404 13685
rect 3399 13574 3451 13626
rect 3463 13574 3515 13626
rect 3527 13574 3579 13626
rect 3591 13574 3643 13626
rect 3655 13574 3707 13626
rect 8298 13574 8350 13626
rect 8362 13574 8414 13626
rect 8426 13574 8478 13626
rect 8490 13574 8542 13626
rect 8554 13574 8606 13626
rect 13197 13574 13249 13626
rect 13261 13574 13313 13626
rect 13325 13574 13377 13626
rect 13389 13574 13441 13626
rect 13453 13574 13505 13626
rect 18096 13574 18148 13626
rect 18160 13574 18212 13626
rect 18224 13574 18276 13626
rect 18288 13574 18340 13626
rect 18352 13574 18404 13626
rect 7840 13515 7892 13524
rect 7840 13481 7849 13515
rect 7849 13481 7883 13515
rect 7883 13481 7892 13515
rect 7840 13472 7892 13481
rect 10508 13472 10560 13524
rect 13084 13515 13136 13524
rect 13084 13481 13093 13515
rect 13093 13481 13127 13515
rect 13127 13481 13136 13515
rect 13084 13472 13136 13481
rect 17408 13515 17460 13524
rect 17408 13481 17417 13515
rect 17417 13481 17451 13515
rect 17451 13481 17460 13515
rect 17408 13472 17460 13481
rect 1492 13311 1544 13320
rect 1492 13277 1501 13311
rect 1501 13277 1535 13311
rect 1535 13277 1544 13311
rect 1492 13268 1544 13277
rect 2228 13379 2280 13388
rect 2228 13345 2237 13379
rect 2237 13345 2271 13379
rect 2271 13345 2280 13379
rect 2228 13336 2280 13345
rect 4896 13268 4948 13320
rect 7380 13311 7432 13320
rect 7380 13277 7389 13311
rect 7389 13277 7423 13311
rect 7423 13277 7432 13311
rect 7380 13268 7432 13277
rect 7840 13268 7892 13320
rect 8484 13268 8536 13320
rect 9588 13268 9640 13320
rect 6920 13132 6972 13184
rect 9864 13268 9916 13320
rect 10416 13311 10468 13320
rect 10416 13277 10425 13311
rect 10425 13277 10459 13311
rect 10459 13277 10468 13311
rect 10416 13268 10468 13277
rect 12532 13404 12584 13456
rect 20168 13447 20220 13456
rect 20168 13413 20177 13447
rect 20177 13413 20211 13447
rect 20211 13413 20220 13447
rect 20168 13404 20220 13413
rect 12164 13379 12216 13388
rect 12164 13345 12173 13379
rect 12173 13345 12207 13379
rect 12207 13345 12216 13379
rect 12164 13336 12216 13345
rect 13912 13336 13964 13388
rect 14372 13379 14424 13388
rect 14372 13345 14381 13379
rect 14381 13345 14415 13379
rect 14415 13345 14424 13379
rect 14372 13336 14424 13345
rect 11980 13268 12032 13320
rect 10600 13200 10652 13252
rect 12532 13311 12584 13320
rect 12532 13277 12541 13311
rect 12541 13277 12575 13311
rect 12575 13277 12584 13311
rect 12532 13268 12584 13277
rect 17408 13268 17460 13320
rect 20352 13311 20404 13320
rect 20352 13277 20361 13311
rect 20361 13277 20395 13311
rect 20395 13277 20404 13311
rect 20352 13268 20404 13277
rect 15384 13200 15436 13252
rect 16580 13200 16632 13252
rect 18972 13200 19024 13252
rect 10324 13132 10376 13184
rect 16028 13132 16080 13184
rect 18052 13132 18104 13184
rect 5848 13030 5900 13082
rect 5912 13030 5964 13082
rect 5976 13030 6028 13082
rect 6040 13030 6092 13082
rect 6104 13030 6156 13082
rect 10747 13030 10799 13082
rect 10811 13030 10863 13082
rect 10875 13030 10927 13082
rect 10939 13030 10991 13082
rect 11003 13030 11055 13082
rect 15646 13030 15698 13082
rect 15710 13030 15762 13082
rect 15774 13030 15826 13082
rect 15838 13030 15890 13082
rect 15902 13030 15954 13082
rect 20545 13030 20597 13082
rect 20609 13030 20661 13082
rect 20673 13030 20725 13082
rect 20737 13030 20789 13082
rect 20801 13030 20853 13082
rect 4896 12971 4948 12980
rect 4896 12937 4905 12971
rect 4905 12937 4939 12971
rect 4939 12937 4948 12971
rect 4896 12928 4948 12937
rect 7380 12928 7432 12980
rect 8668 12928 8720 12980
rect 8484 12903 8536 12912
rect 8484 12869 8493 12903
rect 8493 12869 8527 12903
rect 8527 12869 8536 12903
rect 8484 12860 8536 12869
rect 8944 12860 8996 12912
rect 5172 12835 5224 12844
rect 5172 12801 5181 12835
rect 5181 12801 5215 12835
rect 5215 12801 5224 12835
rect 5172 12792 5224 12801
rect 6920 12792 6972 12844
rect 7840 12835 7892 12844
rect 7840 12801 7849 12835
rect 7849 12801 7883 12835
rect 7883 12801 7892 12835
rect 7840 12792 7892 12801
rect 10232 12835 10284 12844
rect 10232 12801 10241 12835
rect 10241 12801 10275 12835
rect 10275 12801 10284 12835
rect 10232 12792 10284 12801
rect 10416 12792 10468 12844
rect 11980 12971 12032 12980
rect 11980 12937 11989 12971
rect 11989 12937 12023 12971
rect 12023 12937 12032 12971
rect 11980 12928 12032 12937
rect 12532 12928 12584 12980
rect 14556 12928 14608 12980
rect 15108 12928 15160 12980
rect 12164 12835 12216 12844
rect 12164 12801 12182 12835
rect 12182 12801 12216 12835
rect 10324 12767 10376 12776
rect 10324 12733 10333 12767
rect 10333 12733 10367 12767
rect 10367 12733 10376 12767
rect 10324 12724 10376 12733
rect 10600 12767 10652 12776
rect 10600 12733 10609 12767
rect 10609 12733 10643 12767
rect 10643 12733 10652 12767
rect 10600 12724 10652 12733
rect 12164 12792 12216 12801
rect 18052 12792 18104 12844
rect 11060 12656 11112 12708
rect 14372 12656 14424 12708
rect 14648 12656 14700 12708
rect 9864 12588 9916 12640
rect 18420 12631 18472 12640
rect 18420 12597 18429 12631
rect 18429 12597 18463 12631
rect 18463 12597 18472 12631
rect 18420 12588 18472 12597
rect 3399 12486 3451 12538
rect 3463 12486 3515 12538
rect 3527 12486 3579 12538
rect 3591 12486 3643 12538
rect 3655 12486 3707 12538
rect 8298 12486 8350 12538
rect 8362 12486 8414 12538
rect 8426 12486 8478 12538
rect 8490 12486 8542 12538
rect 8554 12486 8606 12538
rect 13197 12486 13249 12538
rect 13261 12486 13313 12538
rect 13325 12486 13377 12538
rect 13389 12486 13441 12538
rect 13453 12486 13505 12538
rect 18096 12486 18148 12538
rect 18160 12486 18212 12538
rect 18224 12486 18276 12538
rect 18288 12486 18340 12538
rect 18352 12486 18404 12538
rect 5172 12384 5224 12436
rect 11060 12384 11112 12436
rect 4988 12223 5040 12232
rect 4988 12189 4997 12223
rect 4997 12189 5031 12223
rect 5031 12189 5040 12223
rect 4988 12180 5040 12189
rect 7380 12180 7432 12232
rect 6184 12087 6236 12096
rect 6184 12053 6193 12087
rect 6193 12053 6227 12087
rect 6227 12053 6236 12087
rect 6184 12044 6236 12053
rect 17224 12427 17276 12436
rect 17224 12393 17233 12427
rect 17233 12393 17267 12427
rect 17267 12393 17276 12427
rect 17224 12384 17276 12393
rect 16396 12316 16448 12368
rect 13912 12248 13964 12300
rect 14648 12291 14700 12300
rect 14648 12257 14657 12291
rect 14657 12257 14691 12291
rect 14691 12257 14700 12291
rect 14648 12248 14700 12257
rect 17592 12316 17644 12368
rect 18420 12180 18472 12232
rect 20352 12223 20404 12232
rect 20352 12189 20361 12223
rect 20361 12189 20395 12223
rect 20395 12189 20404 12223
rect 20352 12180 20404 12189
rect 12440 12112 12492 12164
rect 14648 12112 14700 12164
rect 15108 12112 15160 12164
rect 16396 12155 16448 12164
rect 16396 12121 16405 12155
rect 16405 12121 16439 12155
rect 16439 12121 16448 12155
rect 16396 12112 16448 12121
rect 13636 12044 13688 12096
rect 18880 12044 18932 12096
rect 20168 12087 20220 12096
rect 20168 12053 20177 12087
rect 20177 12053 20211 12087
rect 20211 12053 20220 12087
rect 20168 12044 20220 12053
rect 5848 11942 5900 11994
rect 5912 11942 5964 11994
rect 5976 11942 6028 11994
rect 6040 11942 6092 11994
rect 6104 11942 6156 11994
rect 10747 11942 10799 11994
rect 10811 11942 10863 11994
rect 10875 11942 10927 11994
rect 10939 11942 10991 11994
rect 11003 11942 11055 11994
rect 15646 11942 15698 11994
rect 15710 11942 15762 11994
rect 15774 11942 15826 11994
rect 15838 11942 15890 11994
rect 15902 11942 15954 11994
rect 20545 11942 20597 11994
rect 20609 11942 20661 11994
rect 20673 11942 20725 11994
rect 20737 11942 20789 11994
rect 20801 11942 20853 11994
rect 1492 11704 1544 11756
rect 1768 11679 1820 11688
rect 1768 11645 1777 11679
rect 1777 11645 1811 11679
rect 1811 11645 1820 11679
rect 1768 11636 1820 11645
rect 4988 11840 5040 11892
rect 12440 11840 12492 11892
rect 13820 11840 13872 11892
rect 20352 11883 20404 11892
rect 20352 11849 20361 11883
rect 20361 11849 20395 11883
rect 20395 11849 20404 11883
rect 20352 11840 20404 11849
rect 6184 11704 6236 11756
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 14004 11772 14056 11824
rect 18880 11815 18932 11824
rect 18880 11781 18889 11815
rect 18889 11781 18923 11815
rect 18923 11781 18932 11815
rect 18880 11772 18932 11781
rect 19432 11772 19484 11824
rect 11704 11679 11756 11688
rect 11704 11645 11713 11679
rect 11713 11645 11747 11679
rect 11747 11645 11756 11679
rect 11704 11636 11756 11645
rect 11796 11636 11848 11688
rect 15660 11636 15712 11688
rect 16212 11636 16264 11688
rect 6184 11543 6236 11552
rect 6184 11509 6193 11543
rect 6193 11509 6227 11543
rect 6227 11509 6236 11543
rect 6184 11500 6236 11509
rect 15016 11500 15068 11552
rect 3399 11398 3451 11450
rect 3463 11398 3515 11450
rect 3527 11398 3579 11450
rect 3591 11398 3643 11450
rect 3655 11398 3707 11450
rect 8298 11398 8350 11450
rect 8362 11398 8414 11450
rect 8426 11398 8478 11450
rect 8490 11398 8542 11450
rect 8554 11398 8606 11450
rect 13197 11398 13249 11450
rect 13261 11398 13313 11450
rect 13325 11398 13377 11450
rect 13389 11398 13441 11450
rect 13453 11398 13505 11450
rect 18096 11398 18148 11450
rect 18160 11398 18212 11450
rect 18224 11398 18276 11450
rect 18288 11398 18340 11450
rect 18352 11398 18404 11450
rect 8944 11296 8996 11348
rect 9496 11296 9548 11348
rect 11704 11296 11756 11348
rect 14004 11296 14056 11348
rect 6184 11203 6236 11212
rect 6184 11169 6193 11203
rect 6193 11169 6227 11203
rect 6227 11169 6236 11203
rect 6184 11160 6236 11169
rect 2872 11135 2924 11144
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 6092 11092 6144 11144
rect 9220 11135 9272 11144
rect 9220 11101 9229 11135
rect 9229 11101 9263 11135
rect 9263 11101 9272 11135
rect 9220 11092 9272 11101
rect 7748 11024 7800 11076
rect 8024 11024 8076 11076
rect 9772 11135 9824 11144
rect 9772 11101 9781 11135
rect 9781 11101 9815 11135
rect 9815 11101 9824 11135
rect 9772 11092 9824 11101
rect 9864 11135 9916 11144
rect 9864 11101 9873 11135
rect 9873 11101 9907 11135
rect 9907 11101 9916 11135
rect 9864 11092 9916 11101
rect 11152 11135 11204 11144
rect 11152 11101 11170 11135
rect 11170 11101 11204 11135
rect 9956 11024 10008 11076
rect 11152 11092 11204 11101
rect 11428 11160 11480 11212
rect 12348 11160 12400 11212
rect 15660 11203 15712 11212
rect 15660 11169 15669 11203
rect 15669 11169 15703 11203
rect 15703 11169 15712 11203
rect 15660 11160 15712 11169
rect 17132 11203 17184 11212
rect 17132 11169 17141 11203
rect 17141 11169 17175 11203
rect 17175 11169 17184 11203
rect 17132 11160 17184 11169
rect 14096 11135 14148 11144
rect 14096 11101 14105 11135
rect 14105 11101 14139 11135
rect 14139 11101 14148 11135
rect 14096 11092 14148 11101
rect 2412 10956 2464 11008
rect 6368 10956 6420 11008
rect 7840 10956 7892 11008
rect 15384 10956 15436 11008
rect 5848 10854 5900 10906
rect 5912 10854 5964 10906
rect 5976 10854 6028 10906
rect 6040 10854 6092 10906
rect 6104 10854 6156 10906
rect 10747 10854 10799 10906
rect 10811 10854 10863 10906
rect 10875 10854 10927 10906
rect 10939 10854 10991 10906
rect 11003 10854 11055 10906
rect 15646 10854 15698 10906
rect 15710 10854 15762 10906
rect 15774 10854 15826 10906
rect 15838 10854 15890 10906
rect 15902 10854 15954 10906
rect 20545 10854 20597 10906
rect 20609 10854 20661 10906
rect 20673 10854 20725 10906
rect 20737 10854 20789 10906
rect 20801 10854 20853 10906
rect 3976 10752 4028 10804
rect 8024 10684 8076 10736
rect 9220 10752 9272 10804
rect 9680 10684 9732 10736
rect 2412 10659 2464 10668
rect 2412 10625 2421 10659
rect 2421 10625 2455 10659
rect 2455 10625 2464 10659
rect 2412 10616 2464 10625
rect 6368 10659 6420 10668
rect 6368 10625 6377 10659
rect 6377 10625 6411 10659
rect 6411 10625 6420 10659
rect 6368 10616 6420 10625
rect 7932 10616 7984 10668
rect 11152 10752 11204 10804
rect 11244 10752 11296 10804
rect 11796 10752 11848 10804
rect 14096 10752 14148 10804
rect 17592 10752 17644 10804
rect 19432 10684 19484 10736
rect 11520 10659 11572 10668
rect 7840 10548 7892 10600
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 14464 10616 14516 10668
rect 17132 10616 17184 10668
rect 2320 10412 2372 10464
rect 8116 10455 8168 10464
rect 8116 10421 8125 10455
rect 8125 10421 8159 10455
rect 8159 10421 8168 10455
rect 8116 10412 8168 10421
rect 9128 10548 9180 10600
rect 9772 10548 9824 10600
rect 10968 10548 11020 10600
rect 16396 10548 16448 10600
rect 17408 10548 17460 10600
rect 18604 10591 18656 10600
rect 18604 10557 18613 10591
rect 18613 10557 18647 10591
rect 18647 10557 18656 10591
rect 18604 10548 18656 10557
rect 10048 10412 10100 10464
rect 10508 10455 10560 10464
rect 10508 10421 10517 10455
rect 10517 10421 10551 10455
rect 10551 10421 10560 10455
rect 17224 10480 17276 10532
rect 10508 10412 10560 10421
rect 11888 10412 11940 10464
rect 12164 10412 12216 10464
rect 16580 10412 16632 10464
rect 17500 10412 17552 10464
rect 20352 10455 20404 10464
rect 20352 10421 20361 10455
rect 20361 10421 20395 10455
rect 20395 10421 20404 10455
rect 20352 10412 20404 10421
rect 3399 10310 3451 10362
rect 3463 10310 3515 10362
rect 3527 10310 3579 10362
rect 3591 10310 3643 10362
rect 3655 10310 3707 10362
rect 8298 10310 8350 10362
rect 8362 10310 8414 10362
rect 8426 10310 8478 10362
rect 8490 10310 8542 10362
rect 8554 10310 8606 10362
rect 13197 10310 13249 10362
rect 13261 10310 13313 10362
rect 13325 10310 13377 10362
rect 13389 10310 13441 10362
rect 13453 10310 13505 10362
rect 18096 10310 18148 10362
rect 18160 10310 18212 10362
rect 18224 10310 18276 10362
rect 18288 10310 18340 10362
rect 18352 10310 18404 10362
rect 1768 10208 1820 10260
rect 7932 10251 7984 10260
rect 7932 10217 7941 10251
rect 7941 10217 7975 10251
rect 7975 10217 7984 10251
rect 7932 10208 7984 10217
rect 9128 10251 9180 10260
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 9864 10208 9916 10260
rect 10048 10208 10100 10260
rect 848 10004 900 10056
rect 2320 10047 2372 10056
rect 2320 10013 2329 10047
rect 2329 10013 2363 10047
rect 2363 10013 2372 10047
rect 2320 10004 2372 10013
rect 3976 10004 4028 10056
rect 13176 10183 13228 10192
rect 13176 10149 13185 10183
rect 13185 10149 13219 10183
rect 13219 10149 13228 10183
rect 13176 10140 13228 10149
rect 6276 10072 6328 10124
rect 7840 10004 7892 10056
rect 10232 10072 10284 10124
rect 10508 10004 10560 10056
rect 11244 10072 11296 10124
rect 13084 10072 13136 10124
rect 10968 10047 11020 10056
rect 10968 10013 10977 10047
rect 10977 10013 11011 10047
rect 11011 10013 11020 10047
rect 10968 10004 11020 10013
rect 11428 10047 11480 10056
rect 11428 10013 11437 10047
rect 11437 10013 11471 10047
rect 11471 10013 11480 10047
rect 11428 10004 11480 10013
rect 2964 9936 3016 9988
rect 12164 9936 12216 9988
rect 4528 9868 4580 9920
rect 4712 9868 4764 9920
rect 11520 9868 11572 9920
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 13544 10004 13596 10013
rect 13728 10047 13780 10056
rect 13728 10013 13737 10047
rect 13737 10013 13771 10047
rect 13771 10013 13780 10047
rect 13728 10004 13780 10013
rect 14464 10251 14516 10260
rect 14464 10217 14473 10251
rect 14473 10217 14507 10251
rect 14507 10217 14516 10251
rect 14464 10208 14516 10217
rect 17224 10208 17276 10260
rect 17592 10140 17644 10192
rect 20168 10183 20220 10192
rect 20168 10149 20177 10183
rect 20177 10149 20211 10183
rect 20211 10149 20220 10183
rect 20168 10140 20220 10149
rect 17408 10072 17460 10124
rect 20352 10047 20404 10056
rect 20352 10013 20361 10047
rect 20361 10013 20395 10047
rect 20395 10013 20404 10047
rect 20352 10004 20404 10013
rect 15384 9868 15436 9920
rect 18512 9911 18564 9920
rect 18512 9877 18521 9911
rect 18521 9877 18555 9911
rect 18555 9877 18564 9911
rect 18512 9868 18564 9877
rect 5848 9766 5900 9818
rect 5912 9766 5964 9818
rect 5976 9766 6028 9818
rect 6040 9766 6092 9818
rect 6104 9766 6156 9818
rect 10747 9766 10799 9818
rect 10811 9766 10863 9818
rect 10875 9766 10927 9818
rect 10939 9766 10991 9818
rect 11003 9766 11055 9818
rect 15646 9766 15698 9818
rect 15710 9766 15762 9818
rect 15774 9766 15826 9818
rect 15838 9766 15890 9818
rect 15902 9766 15954 9818
rect 20545 9766 20597 9818
rect 20609 9766 20661 9818
rect 20673 9766 20725 9818
rect 20737 9766 20789 9818
rect 20801 9766 20853 9818
rect 9312 9664 9364 9716
rect 13084 9664 13136 9716
rect 13544 9664 13596 9716
rect 4712 9639 4764 9648
rect 4712 9605 4721 9639
rect 4721 9605 4755 9639
rect 4755 9605 4764 9639
rect 4712 9596 4764 9605
rect 5724 9596 5776 9648
rect 2964 9571 3016 9580
rect 2964 9537 2973 9571
rect 2973 9537 3007 9571
rect 3007 9537 3016 9571
rect 2964 9528 3016 9537
rect 12348 9528 12400 9580
rect 13176 9571 13228 9580
rect 13176 9537 13220 9571
rect 13220 9537 13228 9571
rect 13176 9528 13228 9537
rect 1676 9503 1728 9512
rect 1676 9469 1685 9503
rect 1685 9469 1719 9503
rect 1719 9469 1728 9503
rect 1676 9460 1728 9469
rect 3884 9460 3936 9512
rect 7196 9460 7248 9512
rect 6644 9392 6696 9444
rect 13728 9392 13780 9444
rect 3399 9222 3451 9274
rect 3463 9222 3515 9274
rect 3527 9222 3579 9274
rect 3591 9222 3643 9274
rect 3655 9222 3707 9274
rect 8298 9222 8350 9274
rect 8362 9222 8414 9274
rect 8426 9222 8478 9274
rect 8490 9222 8542 9274
rect 8554 9222 8606 9274
rect 13197 9222 13249 9274
rect 13261 9222 13313 9274
rect 13325 9222 13377 9274
rect 13389 9222 13441 9274
rect 13453 9222 13505 9274
rect 18096 9222 18148 9274
rect 18160 9222 18212 9274
rect 18224 9222 18276 9274
rect 18288 9222 18340 9274
rect 18352 9222 18404 9274
rect 5632 9163 5684 9172
rect 5632 9129 5641 9163
rect 5641 9129 5675 9163
rect 5675 9129 5684 9163
rect 5632 9120 5684 9129
rect 3884 9027 3936 9036
rect 3884 8993 3893 9027
rect 3893 8993 3927 9027
rect 3927 8993 3936 9027
rect 3884 8984 3936 8993
rect 4528 8984 4580 9036
rect 7012 8916 7064 8968
rect 7564 8959 7616 8968
rect 7564 8925 7573 8959
rect 7573 8925 7607 8959
rect 7607 8925 7616 8959
rect 7564 8916 7616 8925
rect 8116 8916 8168 8968
rect 20352 8959 20404 8968
rect 20352 8925 20361 8959
rect 20361 8925 20395 8959
rect 20395 8925 20404 8959
rect 20352 8916 20404 8925
rect 4804 8848 4856 8900
rect 6644 8823 6696 8832
rect 6644 8789 6653 8823
rect 6653 8789 6687 8823
rect 6687 8789 6696 8823
rect 6644 8780 6696 8789
rect 7196 8823 7248 8832
rect 7196 8789 7205 8823
rect 7205 8789 7239 8823
rect 7239 8789 7248 8823
rect 7196 8780 7248 8789
rect 20168 8823 20220 8832
rect 20168 8789 20177 8823
rect 20177 8789 20211 8823
rect 20211 8789 20220 8823
rect 20168 8780 20220 8789
rect 5848 8678 5900 8730
rect 5912 8678 5964 8730
rect 5976 8678 6028 8730
rect 6040 8678 6092 8730
rect 6104 8678 6156 8730
rect 10747 8678 10799 8730
rect 10811 8678 10863 8730
rect 10875 8678 10927 8730
rect 10939 8678 10991 8730
rect 11003 8678 11055 8730
rect 15646 8678 15698 8730
rect 15710 8678 15762 8730
rect 15774 8678 15826 8730
rect 15838 8678 15890 8730
rect 15902 8678 15954 8730
rect 20545 8678 20597 8730
rect 20609 8678 20661 8730
rect 20673 8678 20725 8730
rect 20737 8678 20789 8730
rect 20801 8678 20853 8730
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 8668 8372 8720 8424
rect 8024 8236 8076 8288
rect 9496 8279 9548 8288
rect 9496 8245 9505 8279
rect 9505 8245 9539 8279
rect 9539 8245 9548 8279
rect 9496 8236 9548 8245
rect 11888 8440 11940 8492
rect 12440 8440 12492 8492
rect 12532 8440 12584 8492
rect 16028 8619 16080 8628
rect 16028 8585 16037 8619
rect 16037 8585 16071 8619
rect 16071 8585 16080 8619
rect 16028 8576 16080 8585
rect 16212 8576 16264 8628
rect 20352 8619 20404 8628
rect 20352 8585 20361 8619
rect 20361 8585 20395 8619
rect 20395 8585 20404 8619
rect 20352 8576 20404 8585
rect 15476 8440 15528 8492
rect 18420 8508 18472 8560
rect 18512 8508 18564 8560
rect 19432 8508 19484 8560
rect 17224 8483 17276 8492
rect 17224 8449 17233 8483
rect 17233 8449 17267 8483
rect 17267 8449 17276 8483
rect 17224 8440 17276 8449
rect 17868 8483 17920 8492
rect 17868 8449 17877 8483
rect 17877 8449 17911 8483
rect 17911 8449 17920 8483
rect 17868 8440 17920 8449
rect 17684 8415 17736 8424
rect 17684 8381 17693 8415
rect 17693 8381 17727 8415
rect 17727 8381 17736 8415
rect 17684 8372 17736 8381
rect 18604 8415 18656 8424
rect 18604 8381 18613 8415
rect 18613 8381 18647 8415
rect 18647 8381 18656 8415
rect 18604 8372 18656 8381
rect 16304 8304 16356 8356
rect 17960 8304 18012 8356
rect 10508 8236 10560 8288
rect 11796 8279 11848 8288
rect 11796 8245 11805 8279
rect 11805 8245 11839 8279
rect 11839 8245 11848 8279
rect 11796 8236 11848 8245
rect 11980 8236 12032 8288
rect 14280 8279 14332 8288
rect 14280 8245 14289 8279
rect 14289 8245 14323 8279
rect 14323 8245 14332 8279
rect 14280 8236 14332 8245
rect 17316 8236 17368 8288
rect 18420 8236 18472 8288
rect 3399 8134 3451 8186
rect 3463 8134 3515 8186
rect 3527 8134 3579 8186
rect 3591 8134 3643 8186
rect 3655 8134 3707 8186
rect 8298 8134 8350 8186
rect 8362 8134 8414 8186
rect 8426 8134 8478 8186
rect 8490 8134 8542 8186
rect 8554 8134 8606 8186
rect 13197 8134 13249 8186
rect 13261 8134 13313 8186
rect 13325 8134 13377 8186
rect 13389 8134 13441 8186
rect 13453 8134 13505 8186
rect 18096 8134 18148 8186
rect 18160 8134 18212 8186
rect 18224 8134 18276 8186
rect 18288 8134 18340 8186
rect 18352 8134 18404 8186
rect 3240 8075 3292 8084
rect 3240 8041 3249 8075
rect 3249 8041 3283 8075
rect 3283 8041 3292 8075
rect 3240 8032 3292 8041
rect 8668 8032 8720 8084
rect 9036 8032 9088 8084
rect 6276 7964 6328 8016
rect 2780 7828 2832 7880
rect 2872 7871 2924 7880
rect 2872 7837 2881 7871
rect 2881 7837 2915 7871
rect 2915 7837 2924 7871
rect 2872 7828 2924 7837
rect 4344 7896 4396 7948
rect 2596 7692 2648 7744
rect 4804 7692 4856 7744
rect 7564 7896 7616 7948
rect 8024 7828 8076 7880
rect 6920 7760 6972 7812
rect 8208 7760 8260 7812
rect 7288 7692 7340 7744
rect 9128 7735 9180 7744
rect 9128 7701 9137 7735
rect 9137 7701 9171 7735
rect 9171 7701 9180 7735
rect 9128 7692 9180 7701
rect 10416 7803 10468 7812
rect 10416 7769 10425 7803
rect 10425 7769 10459 7803
rect 10459 7769 10468 7803
rect 10416 7760 10468 7769
rect 10508 7760 10560 7812
rect 11888 8075 11940 8084
rect 11888 8041 11897 8075
rect 11897 8041 11931 8075
rect 11931 8041 11940 8075
rect 11888 8032 11940 8041
rect 18512 8032 18564 8084
rect 11980 7939 12032 7948
rect 11980 7905 11989 7939
rect 11989 7905 12023 7939
rect 12023 7905 12032 7939
rect 11980 7896 12032 7905
rect 14280 7896 14332 7948
rect 16304 7939 16356 7948
rect 16304 7905 16313 7939
rect 16313 7905 16347 7939
rect 16347 7905 16356 7939
rect 16304 7896 16356 7905
rect 16580 7939 16632 7948
rect 16580 7905 16589 7939
rect 16589 7905 16623 7939
rect 16623 7905 16632 7939
rect 16580 7896 16632 7905
rect 18420 7828 18472 7880
rect 12716 7760 12768 7812
rect 14740 7803 14792 7812
rect 14740 7769 14749 7803
rect 14749 7769 14783 7803
rect 14783 7769 14792 7803
rect 14740 7760 14792 7769
rect 12532 7692 12584 7744
rect 13912 7692 13964 7744
rect 14096 7692 14148 7744
rect 18604 7803 18656 7812
rect 18604 7769 18613 7803
rect 18613 7769 18647 7803
rect 18647 7769 18656 7803
rect 18604 7760 18656 7769
rect 5848 7590 5900 7642
rect 5912 7590 5964 7642
rect 5976 7590 6028 7642
rect 6040 7590 6092 7642
rect 6104 7590 6156 7642
rect 10747 7590 10799 7642
rect 10811 7590 10863 7642
rect 10875 7590 10927 7642
rect 10939 7590 10991 7642
rect 11003 7590 11055 7642
rect 15646 7590 15698 7642
rect 15710 7590 15762 7642
rect 15774 7590 15826 7642
rect 15838 7590 15890 7642
rect 15902 7590 15954 7642
rect 20545 7590 20597 7642
rect 20609 7590 20661 7642
rect 20673 7590 20725 7642
rect 20737 7590 20789 7642
rect 20801 7590 20853 7642
rect 4252 7488 4304 7540
rect 4344 7488 4396 7540
rect 7288 7488 7340 7540
rect 10416 7488 10468 7540
rect 3148 7420 3200 7472
rect 5356 7420 5408 7472
rect 9496 7420 9548 7472
rect 2780 7352 2832 7404
rect 2872 7327 2924 7336
rect 2872 7293 2881 7327
rect 2881 7293 2915 7327
rect 2915 7293 2924 7327
rect 2872 7284 2924 7293
rect 3240 7395 3292 7404
rect 3240 7361 3249 7395
rect 3249 7361 3283 7395
rect 3283 7361 3292 7395
rect 3240 7352 3292 7361
rect 7196 7352 7248 7404
rect 8208 7352 8260 7404
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 10508 7352 10560 7404
rect 12440 7531 12492 7540
rect 12440 7497 12449 7531
rect 12449 7497 12483 7531
rect 12483 7497 12492 7531
rect 12440 7488 12492 7497
rect 12716 7488 12768 7540
rect 11796 7463 11848 7472
rect 11796 7429 11805 7463
rect 11805 7429 11839 7463
rect 11839 7429 11848 7463
rect 11796 7420 11848 7429
rect 14096 7488 14148 7540
rect 14740 7488 14792 7540
rect 15476 7531 15528 7540
rect 15476 7497 15485 7531
rect 15485 7497 15519 7531
rect 15519 7497 15528 7531
rect 15476 7488 15528 7497
rect 17224 7488 17276 7540
rect 17684 7531 17736 7540
rect 17684 7497 17693 7531
rect 17693 7497 17727 7531
rect 17727 7497 17736 7531
rect 17684 7488 17736 7497
rect 16580 7352 16632 7404
rect 17316 7395 17368 7404
rect 17316 7361 17325 7395
rect 17325 7361 17359 7395
rect 17359 7361 17368 7395
rect 17316 7352 17368 7361
rect 17960 7395 18012 7404
rect 17960 7361 17969 7395
rect 17969 7361 18003 7395
rect 18003 7361 18012 7395
rect 17960 7352 18012 7361
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 12532 7284 12584 7336
rect 10508 7216 10560 7268
rect 13912 7284 13964 7336
rect 18420 7284 18472 7336
rect 1952 7148 2004 7200
rect 4252 7148 4304 7200
rect 5356 7148 5408 7200
rect 10968 7191 11020 7200
rect 10968 7157 10977 7191
rect 10977 7157 11011 7191
rect 11011 7157 11020 7191
rect 10968 7148 11020 7157
rect 11888 7191 11940 7200
rect 11888 7157 11897 7191
rect 11897 7157 11931 7191
rect 11931 7157 11940 7191
rect 11888 7148 11940 7157
rect 3399 7046 3451 7098
rect 3463 7046 3515 7098
rect 3527 7046 3579 7098
rect 3591 7046 3643 7098
rect 3655 7046 3707 7098
rect 8298 7046 8350 7098
rect 8362 7046 8414 7098
rect 8426 7046 8478 7098
rect 8490 7046 8542 7098
rect 8554 7046 8606 7098
rect 13197 7046 13249 7098
rect 13261 7046 13313 7098
rect 13325 7046 13377 7098
rect 13389 7046 13441 7098
rect 13453 7046 13505 7098
rect 18096 7046 18148 7098
rect 18160 7046 18212 7098
rect 18224 7046 18276 7098
rect 18288 7046 18340 7098
rect 18352 7046 18404 7098
rect 3148 6944 3200 6996
rect 2596 6851 2648 6860
rect 2596 6817 2605 6851
rect 2605 6817 2639 6851
rect 2639 6817 2648 6851
rect 2596 6808 2648 6817
rect 2780 6740 2832 6792
rect 5632 6808 5684 6860
rect 8760 6808 8812 6860
rect 17868 6808 17920 6860
rect 19432 6808 19484 6860
rect 6644 6783 6696 6792
rect 6644 6749 6653 6783
rect 6653 6749 6687 6783
rect 6687 6749 6696 6783
rect 6644 6740 6696 6749
rect 8668 6740 8720 6792
rect 10968 6783 11020 6792
rect 10968 6749 10977 6783
rect 10977 6749 11011 6783
rect 11011 6749 11020 6783
rect 10968 6740 11020 6749
rect 13912 6740 13964 6792
rect 20352 6783 20404 6792
rect 20352 6749 20361 6783
rect 20361 6749 20395 6783
rect 20395 6749 20404 6783
rect 20352 6740 20404 6749
rect 5356 6672 5408 6724
rect 6368 6715 6420 6724
rect 6368 6681 6377 6715
rect 6377 6681 6411 6715
rect 6411 6681 6420 6715
rect 6368 6672 6420 6681
rect 7012 6715 7064 6724
rect 7012 6681 7021 6715
rect 7021 6681 7055 6715
rect 7055 6681 7064 6715
rect 7012 6672 7064 6681
rect 7748 6672 7800 6724
rect 8760 6647 8812 6656
rect 8760 6613 8769 6647
rect 8769 6613 8803 6647
rect 8803 6613 8812 6647
rect 8760 6604 8812 6613
rect 10508 6604 10560 6656
rect 15568 6604 15620 6656
rect 20168 6647 20220 6656
rect 20168 6613 20177 6647
rect 20177 6613 20211 6647
rect 20211 6613 20220 6647
rect 20168 6604 20220 6613
rect 5848 6502 5900 6554
rect 5912 6502 5964 6554
rect 5976 6502 6028 6554
rect 6040 6502 6092 6554
rect 6104 6502 6156 6554
rect 10747 6502 10799 6554
rect 10811 6502 10863 6554
rect 10875 6502 10927 6554
rect 10939 6502 10991 6554
rect 11003 6502 11055 6554
rect 15646 6502 15698 6554
rect 15710 6502 15762 6554
rect 15774 6502 15826 6554
rect 15838 6502 15890 6554
rect 15902 6502 15954 6554
rect 20545 6502 20597 6554
rect 20609 6502 20661 6554
rect 20673 6502 20725 6554
rect 20737 6502 20789 6554
rect 20801 6502 20853 6554
rect 7012 6400 7064 6452
rect 11244 6400 11296 6452
rect 17408 6400 17460 6452
rect 20352 6443 20404 6452
rect 20352 6409 20361 6443
rect 20361 6409 20395 6443
rect 20395 6409 20404 6443
rect 20352 6400 20404 6409
rect 19432 6332 19484 6384
rect 5264 6264 5316 6316
rect 6368 6264 6420 6316
rect 8668 6264 8720 6316
rect 9496 6264 9548 6316
rect 18420 6264 18472 6316
rect 18512 6264 18564 6316
rect 18880 6239 18932 6248
rect 18880 6205 18889 6239
rect 18889 6205 18923 6239
rect 18923 6205 18932 6239
rect 18880 6196 18932 6205
rect 9588 6103 9640 6112
rect 9588 6069 9597 6103
rect 9597 6069 9631 6103
rect 9631 6069 9640 6103
rect 9588 6060 9640 6069
rect 15384 6060 15436 6112
rect 16212 6060 16264 6112
rect 17408 6060 17460 6112
rect 17776 6060 17828 6112
rect 3399 5958 3451 6010
rect 3463 5958 3515 6010
rect 3527 5958 3579 6010
rect 3591 5958 3643 6010
rect 3655 5958 3707 6010
rect 8298 5958 8350 6010
rect 8362 5958 8414 6010
rect 8426 5958 8478 6010
rect 8490 5958 8542 6010
rect 8554 5958 8606 6010
rect 13197 5958 13249 6010
rect 13261 5958 13313 6010
rect 13325 5958 13377 6010
rect 13389 5958 13441 6010
rect 13453 5958 13505 6010
rect 18096 5958 18148 6010
rect 18160 5958 18212 6010
rect 18224 5958 18276 6010
rect 18288 5958 18340 6010
rect 18352 5958 18404 6010
rect 2596 5788 2648 5840
rect 5264 5788 5316 5840
rect 3148 5763 3200 5772
rect 3148 5729 3157 5763
rect 3157 5729 3191 5763
rect 3191 5729 3200 5763
rect 3148 5720 3200 5729
rect 7012 5720 7064 5772
rect 8668 5788 8720 5840
rect 10508 5720 10560 5772
rect 2780 5695 2832 5704
rect 2780 5661 2789 5695
rect 2789 5661 2823 5695
rect 2823 5661 2832 5695
rect 2780 5652 2832 5661
rect 4436 5652 4488 5704
rect 5172 5695 5224 5704
rect 5172 5661 5180 5695
rect 5180 5661 5224 5695
rect 5172 5652 5224 5661
rect 8760 5695 8812 5704
rect 8760 5661 8769 5695
rect 8769 5661 8803 5695
rect 8803 5661 8812 5695
rect 8760 5652 8812 5661
rect 9772 5584 9824 5636
rect 11336 5720 11388 5772
rect 11244 5695 11296 5704
rect 11244 5661 11253 5695
rect 11253 5661 11287 5695
rect 11287 5661 11296 5695
rect 11244 5652 11296 5661
rect 18880 5856 18932 5908
rect 14464 5788 14516 5840
rect 14372 5720 14424 5772
rect 15476 5720 15528 5772
rect 15568 5695 15620 5704
rect 15568 5661 15577 5695
rect 15577 5661 15611 5695
rect 15611 5661 15620 5695
rect 15568 5652 15620 5661
rect 1400 5516 1452 5568
rect 12164 5584 12216 5636
rect 16212 5720 16264 5772
rect 17776 5695 17828 5704
rect 17776 5661 17785 5695
rect 17785 5661 17819 5695
rect 17819 5661 17828 5695
rect 17776 5652 17828 5661
rect 18420 5652 18472 5704
rect 13820 5516 13872 5568
rect 16212 5584 16264 5636
rect 17684 5584 17736 5636
rect 17592 5559 17644 5568
rect 17592 5525 17601 5559
rect 17601 5525 17635 5559
rect 17635 5525 17644 5559
rect 17592 5516 17644 5525
rect 20260 5559 20312 5568
rect 20260 5525 20269 5559
rect 20269 5525 20303 5559
rect 20303 5525 20312 5559
rect 20260 5516 20312 5525
rect 5848 5414 5900 5466
rect 5912 5414 5964 5466
rect 5976 5414 6028 5466
rect 6040 5414 6092 5466
rect 6104 5414 6156 5466
rect 10747 5414 10799 5466
rect 10811 5414 10863 5466
rect 10875 5414 10927 5466
rect 10939 5414 10991 5466
rect 11003 5414 11055 5466
rect 15646 5414 15698 5466
rect 15710 5414 15762 5466
rect 15774 5414 15826 5466
rect 15838 5414 15890 5466
rect 15902 5414 15954 5466
rect 20545 5414 20597 5466
rect 20609 5414 20661 5466
rect 20673 5414 20725 5466
rect 20737 5414 20789 5466
rect 20801 5414 20853 5466
rect 3148 5244 3200 5296
rect 5172 5312 5224 5364
rect 5724 5312 5776 5364
rect 4068 5244 4120 5296
rect 5632 5244 5684 5296
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 2596 5108 2648 5160
rect 3240 4972 3292 5024
rect 4068 5108 4120 5160
rect 5448 5176 5500 5228
rect 7012 5244 7064 5296
rect 8668 5244 8720 5296
rect 5172 5151 5224 5160
rect 5172 5117 5181 5151
rect 5181 5117 5215 5151
rect 5215 5117 5224 5151
rect 5172 5108 5224 5117
rect 6276 5108 6328 5160
rect 14464 5312 14516 5364
rect 16028 5244 16080 5296
rect 18420 5355 18472 5364
rect 18420 5321 18429 5355
rect 18429 5321 18463 5355
rect 18463 5321 18472 5355
rect 18420 5312 18472 5321
rect 19248 5244 19300 5296
rect 19340 5244 19392 5296
rect 9588 5219 9640 5228
rect 9588 5185 9597 5219
rect 9597 5185 9631 5219
rect 9631 5185 9640 5219
rect 9588 5176 9640 5185
rect 12256 5176 12308 5228
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 3792 4972 3844 5024
rect 10508 5040 10560 5092
rect 8208 5015 8260 5024
rect 8208 4981 8217 5015
rect 8217 4981 8251 5015
rect 8251 4981 8260 5015
rect 8208 4972 8260 4981
rect 18788 5151 18840 5160
rect 18788 5117 18797 5151
rect 18797 5117 18831 5151
rect 18831 5117 18840 5151
rect 18788 5108 18840 5117
rect 14096 5040 14148 5092
rect 14372 4972 14424 5024
rect 20076 4972 20128 5024
rect 3399 4870 3451 4922
rect 3463 4870 3515 4922
rect 3527 4870 3579 4922
rect 3591 4870 3643 4922
rect 3655 4870 3707 4922
rect 8298 4870 8350 4922
rect 8362 4870 8414 4922
rect 8426 4870 8478 4922
rect 8490 4870 8542 4922
rect 8554 4870 8606 4922
rect 13197 4870 13249 4922
rect 13261 4870 13313 4922
rect 13325 4870 13377 4922
rect 13389 4870 13441 4922
rect 13453 4870 13505 4922
rect 18096 4870 18148 4922
rect 18160 4870 18212 4922
rect 18224 4870 18276 4922
rect 18288 4870 18340 4922
rect 18352 4870 18404 4922
rect 4436 4811 4488 4820
rect 4436 4777 4445 4811
rect 4445 4777 4479 4811
rect 4479 4777 4488 4811
rect 4436 4768 4488 4777
rect 5172 4768 5224 4820
rect 5448 4768 5500 4820
rect 8668 4768 8720 4820
rect 12256 4811 12308 4820
rect 12256 4777 12265 4811
rect 12265 4777 12299 4811
rect 12299 4777 12308 4811
rect 12256 4768 12308 4777
rect 14096 4811 14148 4820
rect 14096 4777 14105 4811
rect 14105 4777 14139 4811
rect 14139 4777 14148 4811
rect 14096 4768 14148 4777
rect 18788 4768 18840 4820
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 5080 4700 5132 4752
rect 7012 4564 7064 4616
rect 8208 4700 8260 4752
rect 15108 4743 15160 4752
rect 15108 4709 15117 4743
rect 15117 4709 15151 4743
rect 15151 4709 15160 4743
rect 15108 4700 15160 4709
rect 3056 4496 3108 4548
rect 7932 4607 7984 4616
rect 7932 4573 7941 4607
rect 7941 4573 7975 4607
rect 7975 4573 7984 4607
rect 7932 4564 7984 4573
rect 10508 4675 10560 4684
rect 10508 4641 10517 4675
rect 10517 4641 10551 4675
rect 10551 4641 10560 4675
rect 10508 4632 10560 4641
rect 11336 4632 11388 4684
rect 14372 4632 14424 4684
rect 13820 4564 13872 4616
rect 12164 4496 12216 4548
rect 5848 4326 5900 4378
rect 5912 4326 5964 4378
rect 5976 4326 6028 4378
rect 6040 4326 6092 4378
rect 6104 4326 6156 4378
rect 10747 4326 10799 4378
rect 10811 4326 10863 4378
rect 10875 4326 10927 4378
rect 10939 4326 10991 4378
rect 11003 4326 11055 4378
rect 15646 4326 15698 4378
rect 15710 4326 15762 4378
rect 15774 4326 15826 4378
rect 15838 4326 15890 4378
rect 15902 4326 15954 4378
rect 20545 4326 20597 4378
rect 20609 4326 20661 4378
rect 20673 4326 20725 4378
rect 20737 4326 20789 4378
rect 20801 4326 20853 4378
rect 19340 4156 19392 4208
rect 7932 4088 7984 4140
rect 18512 4088 18564 4140
rect 8208 4020 8260 4072
rect 2964 3884 3016 3936
rect 3148 3884 3200 3936
rect 11888 3952 11940 4004
rect 17592 3952 17644 4004
rect 8208 3884 8260 3936
rect 20352 3927 20404 3936
rect 20352 3893 20361 3927
rect 20361 3893 20395 3927
rect 20395 3893 20404 3927
rect 20352 3884 20404 3893
rect 3399 3782 3451 3834
rect 3463 3782 3515 3834
rect 3527 3782 3579 3834
rect 3591 3782 3643 3834
rect 3655 3782 3707 3834
rect 8298 3782 8350 3834
rect 8362 3782 8414 3834
rect 8426 3782 8478 3834
rect 8490 3782 8542 3834
rect 8554 3782 8606 3834
rect 13197 3782 13249 3834
rect 13261 3782 13313 3834
rect 13325 3782 13377 3834
rect 13389 3782 13441 3834
rect 13453 3782 13505 3834
rect 18096 3782 18148 3834
rect 18160 3782 18212 3834
rect 18224 3782 18276 3834
rect 18288 3782 18340 3834
rect 18352 3782 18404 3834
rect 7748 3680 7800 3732
rect 20260 3655 20312 3664
rect 20260 3621 20269 3655
rect 20269 3621 20303 3655
rect 20303 3621 20312 3655
rect 20260 3612 20312 3621
rect 5264 3587 5316 3596
rect 5264 3553 5273 3587
rect 5273 3553 5307 3587
rect 5307 3553 5316 3587
rect 5264 3544 5316 3553
rect 8208 3587 8260 3596
rect 8208 3553 8217 3587
rect 8217 3553 8251 3587
rect 8251 3553 8260 3587
rect 8208 3544 8260 3553
rect 10600 3544 10652 3596
rect 11336 3544 11388 3596
rect 15292 3544 15344 3596
rect 15660 3544 15712 3596
rect 16028 3544 16080 3596
rect 3148 3519 3200 3528
rect 3148 3485 3157 3519
rect 3157 3485 3191 3519
rect 3191 3485 3200 3519
rect 3148 3476 3200 3485
rect 4988 3519 5040 3528
rect 4988 3485 4997 3519
rect 4997 3485 5031 3519
rect 5031 3485 5040 3519
rect 4988 3476 5040 3485
rect 6920 3476 6972 3528
rect 9772 3476 9824 3528
rect 10324 3476 10376 3528
rect 10508 3519 10560 3528
rect 10508 3485 10517 3519
rect 10517 3485 10551 3519
rect 10551 3485 10560 3519
rect 10508 3476 10560 3485
rect 20076 3519 20128 3528
rect 20076 3485 20085 3519
rect 20085 3485 20119 3519
rect 20119 3485 20128 3519
rect 20076 3476 20128 3485
rect 4068 3408 4120 3460
rect 5724 3408 5776 3460
rect 8668 3408 8720 3460
rect 12072 3408 12124 3460
rect 1400 3383 1452 3392
rect 1400 3349 1409 3383
rect 1409 3349 1443 3383
rect 1443 3349 1452 3383
rect 1400 3340 1452 3349
rect 7104 3340 7156 3392
rect 9588 3340 9640 3392
rect 10232 3383 10284 3392
rect 10232 3349 10241 3383
rect 10241 3349 10275 3383
rect 10275 3349 10284 3383
rect 10232 3340 10284 3349
rect 12532 3340 12584 3392
rect 16212 3408 16264 3460
rect 17408 3340 17460 3392
rect 5848 3238 5900 3290
rect 5912 3238 5964 3290
rect 5976 3238 6028 3290
rect 6040 3238 6092 3290
rect 6104 3238 6156 3290
rect 10747 3238 10799 3290
rect 10811 3238 10863 3290
rect 10875 3238 10927 3290
rect 10939 3238 10991 3290
rect 11003 3238 11055 3290
rect 15646 3238 15698 3290
rect 15710 3238 15762 3290
rect 15774 3238 15826 3290
rect 15838 3238 15890 3290
rect 15902 3238 15954 3290
rect 20545 3238 20597 3290
rect 20609 3238 20661 3290
rect 20673 3238 20725 3290
rect 20737 3238 20789 3290
rect 20801 3238 20853 3290
rect 15108 3136 15160 3188
rect 16212 3136 16264 3188
rect 4068 3068 4120 3120
rect 7656 3068 7708 3120
rect 10232 3068 10284 3120
rect 12072 3068 12124 3120
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 4988 3000 5040 3052
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 17132 3000 17184 3052
rect 20352 3043 20404 3052
rect 20352 3009 20361 3043
rect 20361 3009 20395 3043
rect 20395 3009 20404 3043
rect 20352 3000 20404 3009
rect 3056 2932 3108 2984
rect 5264 2932 5316 2984
rect 6276 2932 6328 2984
rect 9496 2932 9548 2984
rect 11888 2932 11940 2984
rect 11336 2864 11388 2916
rect 16028 2932 16080 2984
rect 1492 2839 1544 2848
rect 1492 2805 1501 2839
rect 1501 2805 1535 2839
rect 1535 2805 1544 2839
rect 1492 2796 1544 2805
rect 4436 2796 4488 2848
rect 8668 2796 8720 2848
rect 11244 2796 11296 2848
rect 18972 2796 19024 2848
rect 20168 2839 20220 2848
rect 20168 2805 20177 2839
rect 20177 2805 20211 2839
rect 20211 2805 20220 2839
rect 20168 2796 20220 2805
rect 3399 2694 3451 2746
rect 3463 2694 3515 2746
rect 3527 2694 3579 2746
rect 3591 2694 3643 2746
rect 3655 2694 3707 2746
rect 8298 2694 8350 2746
rect 8362 2694 8414 2746
rect 8426 2694 8478 2746
rect 8490 2694 8542 2746
rect 8554 2694 8606 2746
rect 13197 2694 13249 2746
rect 13261 2694 13313 2746
rect 13325 2694 13377 2746
rect 13389 2694 13441 2746
rect 13453 2694 13505 2746
rect 18096 2694 18148 2746
rect 18160 2694 18212 2746
rect 18224 2694 18276 2746
rect 18288 2694 18340 2746
rect 18352 2694 18404 2746
rect 10324 2592 10376 2644
rect 10600 2524 10652 2576
rect 4988 2456 5040 2508
rect 1400 2388 1452 2440
rect 1952 2431 2004 2440
rect 1952 2397 1961 2431
rect 1961 2397 1995 2431
rect 1995 2397 2004 2431
rect 1952 2388 2004 2397
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 8944 2499 8996 2508
rect 8944 2465 8953 2499
rect 8953 2465 8987 2499
rect 8987 2465 8996 2499
rect 8944 2456 8996 2465
rect 9496 2456 9548 2508
rect 7104 2431 7156 2440
rect 7104 2397 7113 2431
rect 7113 2397 7147 2431
rect 7147 2397 7156 2431
rect 7104 2388 7156 2397
rect 8668 2388 8720 2440
rect 11244 2431 11296 2440
rect 11244 2397 11253 2431
rect 11253 2397 11287 2431
rect 11287 2397 11296 2431
rect 11244 2388 11296 2397
rect 12532 2431 12584 2440
rect 12532 2397 12541 2431
rect 12541 2397 12575 2431
rect 12575 2397 12584 2431
rect 12532 2388 12584 2397
rect 13544 2431 13596 2440
rect 13544 2397 13553 2431
rect 13553 2397 13587 2431
rect 13587 2397 13596 2431
rect 13544 2388 13596 2397
rect 15016 2388 15068 2440
rect 16120 2431 16172 2440
rect 16120 2397 16129 2431
rect 16129 2397 16163 2431
rect 16163 2397 16172 2431
rect 16120 2388 16172 2397
rect 17408 2431 17460 2440
rect 17408 2397 17417 2431
rect 17417 2397 17451 2431
rect 17451 2397 17460 2431
rect 17408 2388 17460 2397
rect 18972 2431 19024 2440
rect 18972 2397 18981 2431
rect 18981 2397 19015 2431
rect 19015 2397 19024 2431
rect 18972 2388 19024 2397
rect 19524 2431 19576 2440
rect 19524 2397 19533 2431
rect 19533 2397 19567 2431
rect 19567 2397 19576 2431
rect 19524 2388 19576 2397
rect 20444 2388 20496 2440
rect 572 2252 624 2304
rect 1860 2252 1912 2304
rect 3148 2252 3200 2304
rect 4804 2320 4856 2372
rect 10508 2320 10560 2372
rect 5264 2252 5316 2304
rect 5724 2252 5776 2304
rect 7012 2252 7064 2304
rect 8300 2252 8352 2304
rect 12164 2252 12216 2304
rect 13452 2252 13504 2304
rect 14740 2252 14792 2304
rect 16028 2252 16080 2304
rect 17316 2252 17368 2304
rect 18604 2252 18656 2304
rect 19892 2252 19944 2304
rect 21180 2252 21232 2304
rect 5848 2150 5900 2202
rect 5912 2150 5964 2202
rect 5976 2150 6028 2202
rect 6040 2150 6092 2202
rect 6104 2150 6156 2202
rect 10747 2150 10799 2202
rect 10811 2150 10863 2202
rect 10875 2150 10927 2202
rect 10939 2150 10991 2202
rect 11003 2150 11055 2202
rect 15646 2150 15698 2202
rect 15710 2150 15762 2202
rect 15774 2150 15826 2202
rect 15838 2150 15890 2202
rect 15902 2150 15954 2202
rect 20545 2150 20597 2202
rect 20609 2150 20661 2202
rect 20673 2150 20725 2202
rect 20737 2150 20789 2202
rect 20801 2150 20853 2202
<< metal2 >>
rect 570 23224 626 24024
rect 1858 23338 1914 24024
rect 1858 23310 1992 23338
rect 1858 23224 1914 23310
rect 584 21690 612 23224
rect 572 21684 624 21690
rect 572 21626 624 21632
rect 1964 21622 1992 23310
rect 3146 23224 3202 24024
rect 4434 23338 4490 24024
rect 4434 23310 4568 23338
rect 4434 23224 4490 23310
rect 3160 21690 3188 23224
rect 3148 21684 3200 21690
rect 3148 21626 3200 21632
rect 4540 21622 4568 23310
rect 5722 23224 5778 24024
rect 7010 23224 7066 24024
rect 8298 23224 8354 24024
rect 9586 23224 9642 24024
rect 10874 23338 10930 24024
rect 10612 23310 10930 23338
rect 5736 21690 5764 23224
rect 5848 21788 6156 21797
rect 5848 21786 5854 21788
rect 5910 21786 5934 21788
rect 5990 21786 6014 21788
rect 6070 21786 6094 21788
rect 6150 21786 6156 21788
rect 5910 21734 5912 21786
rect 6092 21734 6094 21786
rect 5848 21732 5854 21734
rect 5910 21732 5934 21734
rect 5990 21732 6014 21734
rect 6070 21732 6094 21734
rect 6150 21732 6156 21734
rect 5848 21723 6156 21732
rect 7024 21690 7052 23224
rect 8312 21690 8340 23224
rect 5724 21684 5776 21690
rect 5724 21626 5776 21632
rect 7012 21684 7064 21690
rect 7012 21626 7064 21632
rect 8300 21684 8352 21690
rect 8300 21626 8352 21632
rect 9600 21622 9628 23224
rect 10612 21690 10640 23310
rect 10874 23224 10930 23310
rect 12162 23224 12218 24024
rect 13450 23224 13506 24024
rect 14738 23224 14794 24024
rect 16026 23224 16082 24024
rect 17314 23338 17370 24024
rect 17314 23310 17632 23338
rect 17314 23224 17370 23310
rect 10747 21788 11055 21797
rect 10747 21786 10753 21788
rect 10809 21786 10833 21788
rect 10889 21786 10913 21788
rect 10969 21786 10993 21788
rect 11049 21786 11055 21788
rect 10809 21734 10811 21786
rect 10991 21734 10993 21786
rect 10747 21732 10753 21734
rect 10809 21732 10833 21734
rect 10889 21732 10913 21734
rect 10969 21732 10993 21734
rect 11049 21732 11055 21734
rect 10747 21723 11055 21732
rect 10600 21684 10652 21690
rect 10600 21626 10652 21632
rect 12176 21622 12204 23224
rect 13464 21690 13492 23224
rect 14752 21690 14780 23224
rect 15646 21788 15954 21797
rect 15646 21786 15652 21788
rect 15708 21786 15732 21788
rect 15788 21786 15812 21788
rect 15868 21786 15892 21788
rect 15948 21786 15954 21788
rect 15708 21734 15710 21786
rect 15890 21734 15892 21786
rect 15646 21732 15652 21734
rect 15708 21732 15732 21734
rect 15788 21732 15812 21734
rect 15868 21732 15892 21734
rect 15948 21732 15954 21734
rect 15646 21723 15954 21732
rect 16040 21690 16068 23224
rect 17604 21690 17632 23310
rect 18602 23224 18658 24024
rect 19890 23338 19946 24024
rect 19890 23310 20116 23338
rect 19890 23224 19946 23310
rect 18616 21690 18644 23224
rect 20088 21690 20116 23310
rect 21178 23224 21234 24024
rect 20545 21788 20853 21797
rect 20545 21786 20551 21788
rect 20607 21786 20631 21788
rect 20687 21786 20711 21788
rect 20767 21786 20791 21788
rect 20847 21786 20853 21788
rect 20607 21734 20609 21786
rect 20789 21734 20791 21786
rect 20545 21732 20551 21734
rect 20607 21732 20631 21734
rect 20687 21732 20711 21734
rect 20767 21732 20791 21734
rect 20847 21732 20853 21734
rect 20545 21723 20853 21732
rect 13452 21684 13504 21690
rect 13452 21626 13504 21632
rect 14740 21684 14792 21690
rect 14740 21626 14792 21632
rect 16028 21684 16080 21690
rect 16028 21626 16080 21632
rect 17592 21684 17644 21690
rect 17592 21626 17644 21632
rect 18604 21684 18656 21690
rect 18604 21626 18656 21632
rect 20076 21684 20128 21690
rect 20076 21626 20128 21632
rect 1952 21616 2004 21622
rect 1952 21558 2004 21564
rect 4528 21616 4580 21622
rect 4528 21558 4580 21564
rect 9588 21616 9640 21622
rect 9588 21558 9640 21564
rect 12164 21616 12216 21622
rect 12164 21558 12216 21564
rect 19614 21584 19670 21593
rect 1492 21548 1544 21554
rect 1492 21490 1544 21496
rect 3056 21548 3108 21554
rect 3056 21490 3108 21496
rect 3792 21548 3844 21554
rect 3792 21490 3844 21496
rect 4896 21548 4948 21554
rect 4896 21490 4948 21496
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 7196 21548 7248 21554
rect 7196 21490 7248 21496
rect 8852 21548 8904 21554
rect 8852 21490 8904 21496
rect 10048 21548 10100 21554
rect 10048 21490 10100 21496
rect 11612 21548 11664 21554
rect 11612 21490 11664 21496
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 16764 21548 16816 21554
rect 16764 21490 16816 21496
rect 17500 21548 17552 21554
rect 17500 21490 17552 21496
rect 19340 21548 19392 21554
rect 19614 21519 19670 21528
rect 19708 21548 19760 21554
rect 19340 21490 19392 21496
rect 1306 21312 1362 21321
rect 1306 21247 1362 21256
rect 1320 21146 1348 21247
rect 1308 21140 1360 21146
rect 1308 21082 1360 21088
rect 1504 19514 1532 21490
rect 1492 19508 1544 19514
rect 1492 19450 1544 19456
rect 2136 19440 2188 19446
rect 2136 19382 2188 19388
rect 2964 19440 3016 19446
rect 2964 19382 3016 19388
rect 1952 18760 2004 18766
rect 1952 18702 2004 18708
rect 1492 17672 1544 17678
rect 1492 17614 1544 17620
rect 1860 17672 1912 17678
rect 1860 17614 1912 17620
rect 1504 16574 1532 17614
rect 1872 17338 1900 17614
rect 1860 17332 1912 17338
rect 1860 17274 1912 17280
rect 1964 17202 1992 18702
rect 2148 17542 2176 19382
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 2884 18970 2912 19246
rect 2872 18964 2924 18970
rect 2872 18906 2924 18912
rect 2872 17604 2924 17610
rect 2872 17546 2924 17552
rect 2136 17536 2188 17542
rect 2136 17478 2188 17484
rect 1952 17196 2004 17202
rect 1952 17138 2004 17144
rect 1504 16546 1624 16574
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13705 1440 13874
rect 1492 13728 1544 13734
rect 1398 13696 1454 13705
rect 1492 13670 1544 13676
rect 1398 13631 1454 13640
rect 1504 13326 1532 13670
rect 1492 13320 1544 13326
rect 1492 13262 1544 13268
rect 1504 11762 1532 13262
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 848 10056 900 10062
rect 846 10024 848 10033
rect 900 10024 902 10033
rect 846 9959 902 9968
rect 1596 6914 1624 16546
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 15162 1808 15438
rect 2148 15162 2176 17478
rect 2884 17338 2912 17546
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2688 15428 2740 15434
rect 2688 15370 2740 15376
rect 2700 15162 2728 15370
rect 1768 15156 1820 15162
rect 1768 15098 1820 15104
rect 2136 15156 2188 15162
rect 2136 15098 2188 15104
rect 2688 15156 2740 15162
rect 2688 15098 2740 15104
rect 2228 13932 2280 13938
rect 2228 13874 2280 13880
rect 2240 13394 2268 13874
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 1768 11688 1820 11694
rect 1768 11630 1820 11636
rect 1780 10266 1808 11630
rect 2884 11150 2912 16594
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2424 10674 2452 10950
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 2332 10062 2360 10406
rect 2976 10146 3004 19382
rect 3068 15706 3096 21490
rect 3399 21244 3707 21253
rect 3399 21242 3405 21244
rect 3461 21242 3485 21244
rect 3541 21242 3565 21244
rect 3621 21242 3645 21244
rect 3701 21242 3707 21244
rect 3461 21190 3463 21242
rect 3643 21190 3645 21242
rect 3399 21188 3405 21190
rect 3461 21188 3485 21190
rect 3541 21188 3565 21190
rect 3621 21188 3645 21190
rect 3701 21188 3707 21190
rect 3399 21179 3707 21188
rect 3399 20156 3707 20165
rect 3399 20154 3405 20156
rect 3461 20154 3485 20156
rect 3541 20154 3565 20156
rect 3621 20154 3645 20156
rect 3701 20154 3707 20156
rect 3461 20102 3463 20154
rect 3643 20102 3645 20154
rect 3399 20100 3405 20102
rect 3461 20100 3485 20102
rect 3541 20100 3565 20102
rect 3621 20100 3645 20102
rect 3701 20100 3707 20102
rect 3399 20091 3707 20100
rect 3399 19068 3707 19077
rect 3399 19066 3405 19068
rect 3461 19066 3485 19068
rect 3541 19066 3565 19068
rect 3621 19066 3645 19068
rect 3701 19066 3707 19068
rect 3461 19014 3463 19066
rect 3643 19014 3645 19066
rect 3399 19012 3405 19014
rect 3461 19012 3485 19014
rect 3541 19012 3565 19014
rect 3621 19012 3645 19014
rect 3701 19012 3707 19014
rect 3399 19003 3707 19012
rect 3399 17980 3707 17989
rect 3399 17978 3405 17980
rect 3461 17978 3485 17980
rect 3541 17978 3565 17980
rect 3621 17978 3645 17980
rect 3701 17978 3707 17980
rect 3461 17926 3463 17978
rect 3643 17926 3645 17978
rect 3399 17924 3405 17926
rect 3461 17924 3485 17926
rect 3541 17924 3565 17926
rect 3621 17924 3645 17926
rect 3701 17924 3707 17926
rect 3399 17915 3707 17924
rect 3804 17882 3832 21490
rect 4804 20936 4856 20942
rect 4804 20878 4856 20884
rect 3976 20868 4028 20874
rect 3976 20810 4028 20816
rect 3792 17876 3844 17882
rect 3792 17818 3844 17824
rect 3988 17762 4016 20810
rect 4252 20392 4304 20398
rect 4252 20334 4304 20340
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 4080 18766 4108 20198
rect 4264 19854 4292 20334
rect 4816 20058 4844 20878
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 4252 19848 4304 19854
rect 4252 19790 4304 19796
rect 4344 19508 4396 19514
rect 4344 19450 4396 19456
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 4080 18222 4108 18702
rect 4356 18358 4384 19450
rect 4344 18352 4396 18358
rect 4344 18294 4396 18300
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 3804 17734 4016 17762
rect 3516 17536 3568 17542
rect 3516 17478 3568 17484
rect 3528 17202 3556 17478
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 3804 17134 3832 17734
rect 4080 17678 4108 18158
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 3148 16992 3200 16998
rect 3148 16934 3200 16940
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 3160 16590 3188 16934
rect 3252 16658 3280 16934
rect 3399 16892 3707 16901
rect 3399 16890 3405 16892
rect 3461 16890 3485 16892
rect 3541 16890 3565 16892
rect 3621 16890 3645 16892
rect 3701 16890 3707 16892
rect 3461 16838 3463 16890
rect 3643 16838 3645 16890
rect 3399 16836 3405 16838
rect 3461 16836 3485 16838
rect 3541 16836 3565 16838
rect 3621 16836 3645 16838
rect 3701 16836 3707 16838
rect 3399 16827 3707 16836
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3804 16590 3832 17070
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 3792 16584 3844 16590
rect 3792 16526 3844 16532
rect 3399 15804 3707 15813
rect 3399 15802 3405 15804
rect 3461 15802 3485 15804
rect 3541 15802 3565 15804
rect 3621 15802 3645 15804
rect 3701 15802 3707 15804
rect 3461 15750 3463 15802
rect 3643 15750 3645 15802
rect 3399 15748 3405 15750
rect 3461 15748 3485 15750
rect 3541 15748 3565 15750
rect 3621 15748 3645 15750
rect 3701 15748 3707 15750
rect 3399 15739 3707 15748
rect 3988 15706 4016 16934
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 3976 15700 4028 15706
rect 3976 15642 4028 15648
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 3056 14952 3108 14958
rect 3056 14894 3108 14900
rect 2884 10118 3004 10146
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1412 6886 1624 6914
rect 1412 5574 1440 6886
rect 1400 5568 1452 5574
rect 1400 5510 1452 5516
rect 1412 5234 1440 5510
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 1412 2446 1440 3334
rect 1688 3058 1716 9454
rect 2884 7970 2912 10118
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2976 9586 3004 9930
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2884 7942 3004 7970
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 572 2304 624 2310
rect 1504 2281 1532 2790
rect 1964 2446 1992 7142
rect 2608 6866 2636 7686
rect 2792 7410 2820 7822
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2884 7342 2912 7822
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2596 6860 2648 6866
rect 2596 6802 2648 6808
rect 2608 5846 2636 6802
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2596 5840 2648 5846
rect 2596 5782 2648 5788
rect 2608 5166 2636 5782
rect 2792 5710 2820 6734
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 2976 3942 3004 7942
rect 3068 4554 3096 14894
rect 3252 8090 3280 15506
rect 3344 15026 3372 15642
rect 3988 15502 4016 15642
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3516 15360 3568 15366
rect 3516 15302 3568 15308
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 3528 15026 3556 15302
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3399 14716 3707 14725
rect 3399 14714 3405 14716
rect 3461 14714 3485 14716
rect 3541 14714 3565 14716
rect 3621 14714 3645 14716
rect 3701 14714 3707 14716
rect 3461 14662 3463 14714
rect 3643 14662 3645 14714
rect 3399 14660 3405 14662
rect 3461 14660 3485 14662
rect 3541 14660 3565 14662
rect 3621 14660 3645 14662
rect 3701 14660 3707 14662
rect 3399 14651 3707 14660
rect 3988 13870 4016 15302
rect 4908 15162 4936 21490
rect 5080 20800 5132 20806
rect 5080 20742 5132 20748
rect 5092 20398 5120 20742
rect 5080 20392 5132 20398
rect 5080 20334 5132 20340
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 5368 19446 5396 20198
rect 5356 19440 5408 19446
rect 5356 19382 5408 19388
rect 5172 19168 5224 19174
rect 5172 19110 5224 19116
rect 5184 18766 5212 19110
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 5000 15502 5028 16390
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 5184 14618 5212 14894
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 3399 13628 3707 13637
rect 3399 13626 3405 13628
rect 3461 13626 3485 13628
rect 3541 13626 3565 13628
rect 3621 13626 3645 13628
rect 3701 13626 3707 13628
rect 3461 13574 3463 13626
rect 3643 13574 3645 13626
rect 3399 13572 3405 13574
rect 3461 13572 3485 13574
rect 3541 13572 3565 13574
rect 3621 13572 3645 13574
rect 3701 13572 3707 13574
rect 3399 13563 3707 13572
rect 3399 12540 3707 12549
rect 3399 12538 3405 12540
rect 3461 12538 3485 12540
rect 3541 12538 3565 12540
rect 3621 12538 3645 12540
rect 3701 12538 3707 12540
rect 3461 12486 3463 12538
rect 3643 12486 3645 12538
rect 3399 12484 3405 12486
rect 3461 12484 3485 12486
rect 3541 12484 3565 12486
rect 3621 12484 3645 12486
rect 3701 12484 3707 12486
rect 3399 12475 3707 12484
rect 3399 11452 3707 11461
rect 3399 11450 3405 11452
rect 3461 11450 3485 11452
rect 3541 11450 3565 11452
rect 3621 11450 3645 11452
rect 3701 11450 3707 11452
rect 3461 11398 3463 11450
rect 3643 11398 3645 11450
rect 3399 11396 3405 11398
rect 3461 11396 3485 11398
rect 3541 11396 3565 11398
rect 3621 11396 3645 11398
rect 3701 11396 3707 11398
rect 3399 11387 3707 11396
rect 3988 10810 4016 13806
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4908 12986 4936 13262
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 5000 12434 5028 14350
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5184 12442 5212 12786
rect 4908 12406 5028 12434
rect 5172 12436 5224 12442
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3399 10364 3707 10373
rect 3399 10362 3405 10364
rect 3461 10362 3485 10364
rect 3541 10362 3565 10364
rect 3621 10362 3645 10364
rect 3701 10362 3707 10364
rect 3461 10310 3463 10362
rect 3643 10310 3645 10362
rect 3399 10308 3405 10310
rect 3461 10308 3485 10310
rect 3541 10308 3565 10310
rect 3621 10308 3645 10310
rect 3701 10308 3707 10310
rect 3399 10299 3707 10308
rect 3988 10062 4016 10746
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3399 9276 3707 9285
rect 3399 9274 3405 9276
rect 3461 9274 3485 9276
rect 3541 9274 3565 9276
rect 3621 9274 3645 9276
rect 3701 9274 3707 9276
rect 3461 9222 3463 9274
rect 3643 9222 3645 9274
rect 3399 9220 3405 9222
rect 3461 9220 3485 9222
rect 3541 9220 3565 9222
rect 3621 9220 3645 9222
rect 3701 9220 3707 9222
rect 3399 9211 3707 9220
rect 3896 9042 3924 9454
rect 4540 9042 4568 9862
rect 4724 9654 4752 9862
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 3884 9036 3936 9042
rect 3884 8978 3936 8984
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4804 8900 4856 8906
rect 4804 8842 4856 8848
rect 3399 8188 3707 8197
rect 3399 8186 3405 8188
rect 3461 8186 3485 8188
rect 3541 8186 3565 8188
rect 3621 8186 3645 8188
rect 3701 8186 3707 8188
rect 3461 8134 3463 8186
rect 3643 8134 3645 8186
rect 3399 8132 3405 8134
rect 3461 8132 3485 8134
rect 3541 8132 3565 8134
rect 3621 8132 3645 8134
rect 3701 8132 3707 8134
rect 3399 8123 3707 8132
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3160 7002 3188 7414
rect 3252 7410 3280 8026
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4356 7546 4384 7890
rect 4816 7750 4844 8842
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 4264 7206 4292 7482
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 3399 7100 3707 7109
rect 3399 7098 3405 7100
rect 3461 7098 3485 7100
rect 3541 7098 3565 7100
rect 3621 7098 3645 7100
rect 3701 7098 3707 7100
rect 3461 7046 3463 7098
rect 3643 7046 3645 7098
rect 3399 7044 3405 7046
rect 3461 7044 3485 7046
rect 3541 7044 3565 7046
rect 3621 7044 3645 7046
rect 3701 7044 3707 7046
rect 3399 7035 3707 7044
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3399 6012 3707 6021
rect 3399 6010 3405 6012
rect 3461 6010 3485 6012
rect 3541 6010 3565 6012
rect 3621 6010 3645 6012
rect 3701 6010 3707 6012
rect 3461 5958 3463 6010
rect 3643 5958 3645 6010
rect 3399 5956 3405 5958
rect 3461 5956 3485 5958
rect 3541 5956 3565 5958
rect 3621 5956 3645 5958
rect 3701 5956 3707 5958
rect 3399 5947 3707 5956
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 3160 5302 3188 5714
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 3148 5296 3200 5302
rect 3148 5238 3200 5244
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 4080 5166 4108 5238
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 3068 2990 3096 4490
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 3160 3534 3188 3878
rect 3148 3528 3200 3534
rect 3148 3470 3200 3476
rect 3056 2984 3108 2990
rect 3056 2926 3108 2932
rect 3252 2446 3280 4966
rect 3399 4924 3707 4933
rect 3399 4922 3405 4924
rect 3461 4922 3485 4924
rect 3541 4922 3565 4924
rect 3621 4922 3645 4924
rect 3701 4922 3707 4924
rect 3461 4870 3463 4922
rect 3643 4870 3645 4922
rect 3399 4868 3405 4870
rect 3461 4868 3485 4870
rect 3541 4868 3565 4870
rect 3621 4868 3645 4870
rect 3701 4868 3707 4870
rect 3399 4859 3707 4868
rect 3804 4622 3832 4966
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3399 3836 3707 3845
rect 3399 3834 3405 3836
rect 3461 3834 3485 3836
rect 3541 3834 3565 3836
rect 3621 3834 3645 3836
rect 3701 3834 3707 3836
rect 3461 3782 3463 3834
rect 3643 3782 3645 3834
rect 3399 3780 3405 3782
rect 3461 3780 3485 3782
rect 3541 3780 3565 3782
rect 3621 3780 3645 3782
rect 3701 3780 3707 3782
rect 3399 3771 3707 3780
rect 4080 3466 4108 5102
rect 4448 4826 4476 5646
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4080 3126 4108 3402
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 4436 2848 4488 2854
rect 4436 2790 4488 2796
rect 3399 2748 3707 2757
rect 3399 2746 3405 2748
rect 3461 2746 3485 2748
rect 3541 2746 3565 2748
rect 3621 2746 3645 2748
rect 3701 2746 3707 2748
rect 3461 2694 3463 2746
rect 3643 2694 3645 2746
rect 3399 2692 3405 2694
rect 3461 2692 3485 2694
rect 3541 2692 3565 2694
rect 3621 2692 3645 2694
rect 3701 2692 3707 2694
rect 3399 2683 3707 2692
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 1860 2304 1912 2310
rect 572 2246 624 2252
rect 1490 2272 1546 2281
rect 584 800 612 2246
rect 1860 2246 1912 2252
rect 3148 2304 3200 2310
rect 3148 2246 3200 2252
rect 1490 2207 1546 2216
rect 1872 800 1900 2246
rect 3160 800 3188 2246
rect 4448 800 4476 2790
rect 4816 2378 4844 7686
rect 4908 6225 4936 12406
rect 5172 12378 5224 12384
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 5000 11898 5028 12174
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 5644 9178 5672 21490
rect 6736 20868 6788 20874
rect 6736 20810 6788 20816
rect 5848 20700 6156 20709
rect 5848 20698 5854 20700
rect 5910 20698 5934 20700
rect 5990 20698 6014 20700
rect 6070 20698 6094 20700
rect 6150 20698 6156 20700
rect 5910 20646 5912 20698
rect 6092 20646 6094 20698
rect 5848 20644 5854 20646
rect 5910 20644 5934 20646
rect 5990 20644 6014 20646
rect 6070 20644 6094 20646
rect 6150 20644 6156 20646
rect 5848 20635 6156 20644
rect 6748 20534 6776 20810
rect 6736 20528 6788 20534
rect 6736 20470 6788 20476
rect 5848 19612 6156 19621
rect 5848 19610 5854 19612
rect 5910 19610 5934 19612
rect 5990 19610 6014 19612
rect 6070 19610 6094 19612
rect 6150 19610 6156 19612
rect 5910 19558 5912 19610
rect 6092 19558 6094 19610
rect 5848 19556 5854 19558
rect 5910 19556 5934 19558
rect 5990 19556 6014 19558
rect 6070 19556 6094 19558
rect 6150 19556 6156 19558
rect 5848 19547 6156 19556
rect 6748 19514 6776 20470
rect 7012 20392 7064 20398
rect 7012 20334 7064 20340
rect 6736 19508 6788 19514
rect 6736 19450 6788 19456
rect 6748 18698 6776 19450
rect 5724 18692 5776 18698
rect 5724 18634 5776 18640
rect 6736 18692 6788 18698
rect 6736 18634 6788 18640
rect 5736 18426 5764 18634
rect 5848 18524 6156 18533
rect 5848 18522 5854 18524
rect 5910 18522 5934 18524
rect 5990 18522 6014 18524
rect 6070 18522 6094 18524
rect 6150 18522 6156 18524
rect 5910 18470 5912 18522
rect 6092 18470 6094 18522
rect 5848 18468 5854 18470
rect 5910 18468 5934 18470
rect 5990 18468 6014 18470
rect 6070 18468 6094 18470
rect 6150 18468 6156 18470
rect 5848 18459 6156 18468
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 6748 18358 6776 18634
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6736 18352 6788 18358
rect 6736 18294 6788 18300
rect 6748 17542 6776 18294
rect 6932 17746 6960 18566
rect 7024 18222 7052 20334
rect 7012 18216 7064 18222
rect 7012 18158 7064 18164
rect 7024 17882 7052 18158
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 6920 17740 6972 17746
rect 6920 17682 6972 17688
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 5848 17436 6156 17445
rect 5848 17434 5854 17436
rect 5910 17434 5934 17436
rect 5990 17434 6014 17436
rect 6070 17434 6094 17436
rect 6150 17434 6156 17436
rect 5910 17382 5912 17434
rect 6092 17382 6094 17434
rect 5848 17380 5854 17382
rect 5910 17380 5934 17382
rect 5990 17380 6014 17382
rect 6070 17380 6094 17382
rect 6150 17380 6156 17382
rect 5848 17371 6156 17380
rect 5848 16348 6156 16357
rect 5848 16346 5854 16348
rect 5910 16346 5934 16348
rect 5990 16346 6014 16348
rect 6070 16346 6094 16348
rect 6150 16346 6156 16348
rect 5910 16294 5912 16346
rect 6092 16294 6094 16346
rect 5848 16292 5854 16294
rect 5910 16292 5934 16294
rect 5990 16292 6014 16294
rect 6070 16292 6094 16294
rect 6150 16292 6156 16294
rect 5848 16283 6156 16292
rect 6184 16108 6236 16114
rect 6184 16050 6236 16056
rect 5848 15260 6156 15269
rect 5848 15258 5854 15260
rect 5910 15258 5934 15260
rect 5990 15258 6014 15260
rect 6070 15258 6094 15260
rect 6150 15258 6156 15260
rect 5910 15206 5912 15258
rect 6092 15206 6094 15258
rect 5848 15204 5854 15206
rect 5910 15204 5934 15206
rect 5990 15204 6014 15206
rect 6070 15204 6094 15206
rect 6150 15204 6156 15206
rect 5848 15195 6156 15204
rect 6196 15162 6224 16050
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 6380 15026 6408 15846
rect 6368 15020 6420 15026
rect 6368 14962 6420 14968
rect 5848 14172 6156 14181
rect 5848 14170 5854 14172
rect 5910 14170 5934 14172
rect 5990 14170 6014 14172
rect 6070 14170 6094 14172
rect 6150 14170 6156 14172
rect 5910 14118 5912 14170
rect 6092 14118 6094 14170
rect 5848 14116 5854 14118
rect 5910 14116 5934 14118
rect 5990 14116 6014 14118
rect 6070 14116 6094 14118
rect 6150 14116 6156 14118
rect 5848 14107 6156 14116
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 5848 13084 6156 13093
rect 5848 13082 5854 13084
rect 5910 13082 5934 13084
rect 5990 13082 6014 13084
rect 6070 13082 6094 13084
rect 6150 13082 6156 13084
rect 5910 13030 5912 13082
rect 6092 13030 6094 13082
rect 5848 13028 5854 13030
rect 5910 13028 5934 13030
rect 5990 13028 6014 13030
rect 6070 13028 6094 13030
rect 6150 13028 6156 13030
rect 5848 13019 6156 13028
rect 6932 12850 6960 13126
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6932 12434 6960 12786
rect 6932 12406 7052 12434
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 5848 11996 6156 12005
rect 5848 11994 5854 11996
rect 5910 11994 5934 11996
rect 5990 11994 6014 11996
rect 6070 11994 6094 11996
rect 6150 11994 6156 11996
rect 5910 11942 5912 11994
rect 6092 11942 6094 11994
rect 5848 11940 5854 11942
rect 5910 11940 5934 11942
rect 5990 11940 6014 11942
rect 6070 11940 6094 11942
rect 6150 11940 6156 11942
rect 5848 11931 6156 11940
rect 6196 11762 6224 12038
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6196 11642 6224 11698
rect 6104 11614 6224 11642
rect 6104 11150 6132 11614
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6196 11218 6224 11494
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 5848 10908 6156 10917
rect 5848 10906 5854 10908
rect 5910 10906 5934 10908
rect 5990 10906 6014 10908
rect 6070 10906 6094 10908
rect 6150 10906 6156 10908
rect 5910 10854 5912 10906
rect 6092 10854 6094 10906
rect 5848 10852 5854 10854
rect 5910 10852 5934 10854
rect 5990 10852 6014 10854
rect 6070 10852 6094 10854
rect 6150 10852 6156 10854
rect 5848 10843 6156 10852
rect 6380 10674 6408 10950
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 5848 9820 6156 9829
rect 5848 9818 5854 9820
rect 5910 9818 5934 9820
rect 5990 9818 6014 9820
rect 6070 9818 6094 9820
rect 6150 9818 6156 9820
rect 5910 9766 5912 9818
rect 6092 9766 6094 9818
rect 5848 9764 5854 9766
rect 5910 9764 5934 9766
rect 5990 9764 6014 9766
rect 6070 9764 6094 9766
rect 6150 9764 6156 9766
rect 5848 9755 6156 9764
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5368 7206 5396 7414
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5368 6730 5396 7142
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5356 6724 5408 6730
rect 5356 6666 5408 6672
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 4894 6216 4950 6225
rect 4894 6151 4950 6160
rect 5276 5846 5304 6258
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 5184 5370 5212 5646
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5184 5250 5212 5306
rect 5092 5222 5212 5250
rect 5092 4758 5120 5222
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 5184 4826 5212 5102
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5080 4752 5132 4758
rect 5080 4694 5132 4700
rect 5276 3602 5304 5782
rect 5368 5250 5396 6666
rect 5644 5302 5672 6802
rect 5736 5370 5764 9590
rect 5848 8732 6156 8741
rect 5848 8730 5854 8732
rect 5910 8730 5934 8732
rect 5990 8730 6014 8732
rect 6070 8730 6094 8732
rect 6150 8730 6156 8732
rect 5910 8678 5912 8730
rect 6092 8678 6094 8730
rect 5848 8676 5854 8678
rect 5910 8676 5934 8678
rect 5990 8676 6014 8678
rect 6070 8676 6094 8678
rect 6150 8676 6156 8678
rect 5848 8667 6156 8676
rect 6288 8022 6316 10066
rect 6644 9444 6696 9450
rect 6644 9386 6696 9392
rect 6656 8838 6684 9386
rect 7024 8974 7052 12406
rect 7208 9518 7236 21490
rect 8298 21244 8606 21253
rect 8298 21242 8304 21244
rect 8360 21242 8384 21244
rect 8440 21242 8464 21244
rect 8520 21242 8544 21244
rect 8600 21242 8606 21244
rect 8360 21190 8362 21242
rect 8542 21190 8544 21242
rect 8298 21188 8304 21190
rect 8360 21188 8384 21190
rect 8440 21188 8464 21190
rect 8520 21188 8544 21190
rect 8600 21188 8606 21190
rect 8298 21179 8606 21188
rect 7288 20936 7340 20942
rect 7288 20878 7340 20884
rect 8208 20936 8260 20942
rect 8208 20878 8260 20884
rect 7300 20398 7328 20878
rect 7840 20868 7892 20874
rect 7840 20810 7892 20816
rect 7288 20392 7340 20398
rect 7288 20334 7340 20340
rect 7656 20392 7708 20398
rect 7656 20334 7708 20340
rect 7668 20058 7696 20334
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7852 19378 7880 20810
rect 8220 19802 8248 20878
rect 8298 20156 8606 20165
rect 8298 20154 8304 20156
rect 8360 20154 8384 20156
rect 8440 20154 8464 20156
rect 8520 20154 8544 20156
rect 8600 20154 8606 20156
rect 8360 20102 8362 20154
rect 8542 20102 8544 20154
rect 8298 20100 8304 20102
rect 8360 20100 8384 20102
rect 8440 20100 8464 20102
rect 8520 20100 8544 20102
rect 8600 20100 8606 20102
rect 8298 20091 8606 20100
rect 8392 19848 8444 19854
rect 8220 19796 8392 19802
rect 8220 19790 8444 19796
rect 8220 19774 8432 19790
rect 8864 19394 8892 21490
rect 8944 21004 8996 21010
rect 8944 20946 8996 20952
rect 8956 20058 8984 20946
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 9312 20868 9364 20874
rect 9312 20810 9364 20816
rect 9036 20800 9088 20806
rect 9036 20742 9088 20748
rect 9048 20534 9076 20742
rect 9036 20528 9088 20534
rect 9036 20470 9088 20476
rect 8944 20052 8996 20058
rect 8944 19994 8996 20000
rect 8944 19780 8996 19786
rect 9048 19768 9076 20470
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 9140 19854 9168 20198
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 8996 19740 9076 19768
rect 8944 19722 8996 19728
rect 9048 19446 9076 19740
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 8772 19366 8892 19394
rect 9036 19440 9088 19446
rect 9036 19382 9088 19388
rect 8036 18834 8064 19314
rect 8298 19068 8606 19077
rect 8298 19066 8304 19068
rect 8360 19066 8384 19068
rect 8440 19066 8464 19068
rect 8520 19066 8544 19068
rect 8600 19066 8606 19068
rect 8360 19014 8362 19066
rect 8542 19014 8544 19066
rect 8298 19012 8304 19014
rect 8360 19012 8384 19014
rect 8440 19012 8464 19014
rect 8520 19012 8544 19014
rect 8600 19012 8606 19014
rect 8298 19003 8606 19012
rect 8024 18828 8076 18834
rect 8024 18770 8076 18776
rect 8036 18222 8064 18770
rect 7840 18216 7892 18222
rect 7840 18158 7892 18164
rect 8024 18216 8076 18222
rect 8024 18158 8076 18164
rect 7852 17882 7880 18158
rect 8298 17980 8606 17989
rect 8298 17978 8304 17980
rect 8360 17978 8384 17980
rect 8440 17978 8464 17980
rect 8520 17978 8544 17980
rect 8600 17978 8606 17980
rect 8360 17926 8362 17978
rect 8542 17926 8544 17978
rect 8298 17924 8304 17926
rect 8360 17924 8384 17926
rect 8440 17924 8464 17926
rect 8520 17924 8544 17926
rect 8600 17924 8606 17926
rect 8298 17915 8606 17924
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 8298 16892 8606 16901
rect 8298 16890 8304 16892
rect 8360 16890 8384 16892
rect 8440 16890 8464 16892
rect 8520 16890 8544 16892
rect 8600 16890 8606 16892
rect 8360 16838 8362 16890
rect 8542 16838 8544 16890
rect 8298 16836 8304 16838
rect 8360 16836 8384 16838
rect 8440 16836 8464 16838
rect 8520 16836 8544 16838
rect 8600 16836 8606 16838
rect 8298 16827 8606 16836
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 7840 16176 7892 16182
rect 7760 16124 7840 16130
rect 7760 16118 7892 16124
rect 7760 16102 7880 16118
rect 7760 15502 7788 16102
rect 8036 16046 8064 16526
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7760 15366 7788 15438
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 7380 15156 7432 15162
rect 7380 15098 7432 15104
rect 7392 13326 7420 15098
rect 7760 15026 7788 15302
rect 8036 15162 8064 15982
rect 8298 15804 8606 15813
rect 8298 15802 8304 15804
rect 8360 15802 8384 15804
rect 8440 15802 8464 15804
rect 8520 15802 8544 15804
rect 8600 15802 8606 15804
rect 8360 15750 8362 15802
rect 8542 15750 8544 15802
rect 8298 15748 8304 15750
rect 8360 15748 8384 15750
rect 8440 15748 8464 15750
rect 8520 15748 8544 15750
rect 8600 15748 8606 15750
rect 8298 15739 8606 15748
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 8404 15162 8432 15438
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 8392 15156 8444 15162
rect 8392 15098 8444 15104
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7392 12986 7420 13262
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7392 12238 7420 12922
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7760 11082 7788 14962
rect 8298 14716 8606 14725
rect 8298 14714 8304 14716
rect 8360 14714 8384 14716
rect 8440 14714 8464 14716
rect 8520 14714 8544 14716
rect 8600 14714 8606 14716
rect 8360 14662 8362 14714
rect 8542 14662 8544 14714
rect 8298 14660 8304 14662
rect 8360 14660 8384 14662
rect 8440 14660 8464 14662
rect 8520 14660 8544 14662
rect 8600 14660 8606 14662
rect 8298 14651 8606 14660
rect 8680 14006 8708 15302
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7852 13530 7880 13806
rect 8298 13628 8606 13637
rect 8298 13626 8304 13628
rect 8360 13626 8384 13628
rect 8440 13626 8464 13628
rect 8520 13626 8544 13628
rect 8600 13626 8606 13628
rect 8360 13574 8362 13626
rect 8542 13574 8544 13626
rect 8298 13572 8304 13574
rect 8360 13572 8384 13574
rect 8440 13572 8464 13574
rect 8520 13572 8544 13574
rect 8600 13572 8606 13574
rect 8298 13563 8606 13572
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 7852 12850 7880 13262
rect 8496 12918 8524 13262
rect 8680 12986 8708 13942
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 8298 12540 8606 12549
rect 8298 12538 8304 12540
rect 8360 12538 8384 12540
rect 8440 12538 8464 12540
rect 8520 12538 8544 12540
rect 8600 12538 8606 12540
rect 8360 12486 8362 12538
rect 8542 12486 8544 12538
rect 8298 12484 8304 12486
rect 8360 12484 8384 12486
rect 8440 12484 8464 12486
rect 8520 12484 8544 12486
rect 8600 12484 8606 12486
rect 8298 12475 8606 12484
rect 8298 11452 8606 11461
rect 8298 11450 8304 11452
rect 8360 11450 8384 11452
rect 8440 11450 8464 11452
rect 8520 11450 8544 11452
rect 8600 11450 8606 11452
rect 8360 11398 8362 11450
rect 8542 11398 8544 11450
rect 8298 11396 8304 11398
rect 8360 11396 8384 11398
rect 8440 11396 8464 11398
rect 8520 11396 8544 11398
rect 8600 11396 8606 11398
rect 8298 11387 8606 11396
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 7840 11008 7892 11014
rect 7840 10950 7892 10956
rect 7852 10606 7880 10950
rect 8036 10742 8064 11018
rect 8024 10736 8076 10742
rect 8024 10678 8076 10684
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 7852 10062 7880 10542
rect 7944 10266 7972 10610
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 6276 8016 6328 8022
rect 6276 7958 6328 7964
rect 5848 7644 6156 7653
rect 5848 7642 5854 7644
rect 5910 7642 5934 7644
rect 5990 7642 6014 7644
rect 6070 7642 6094 7644
rect 6150 7642 6156 7644
rect 5910 7590 5912 7642
rect 6092 7590 6094 7642
rect 5848 7588 5854 7590
rect 5910 7588 5934 7590
rect 5990 7588 6014 7590
rect 6070 7588 6094 7590
rect 6150 7588 6156 7590
rect 5848 7579 6156 7588
rect 5848 6556 6156 6565
rect 5848 6554 5854 6556
rect 5910 6554 5934 6556
rect 5990 6554 6014 6556
rect 6070 6554 6094 6556
rect 6150 6554 6156 6556
rect 5910 6502 5912 6554
rect 6092 6502 6094 6554
rect 5848 6500 5854 6502
rect 5910 6500 5934 6502
rect 5990 6500 6014 6502
rect 6070 6500 6094 6502
rect 6150 6500 6156 6502
rect 5848 6491 6156 6500
rect 5848 5468 6156 5477
rect 5848 5466 5854 5468
rect 5910 5466 5934 5468
rect 5990 5466 6014 5468
rect 6070 5466 6094 5468
rect 6150 5466 6156 5468
rect 5910 5414 5912 5466
rect 6092 5414 6094 5466
rect 5848 5412 5854 5414
rect 5910 5412 5934 5414
rect 5990 5412 6014 5414
rect 6070 5412 6094 5414
rect 6150 5412 6156 5414
rect 5848 5403 6156 5412
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5632 5296 5684 5302
rect 5368 5234 5488 5250
rect 5632 5238 5684 5244
rect 5368 5228 5500 5234
rect 5368 5222 5448 5228
rect 5448 5170 5500 5176
rect 5460 4826 5488 5170
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 5000 3058 5028 3470
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 5000 2514 5028 2994
rect 5276 2990 5304 3538
rect 5736 3466 5764 5306
rect 6288 5166 6316 7958
rect 6656 6798 6684 8774
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6368 6724 6420 6730
rect 6368 6666 6420 6672
rect 6380 6322 6408 6666
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6276 5160 6328 5166
rect 6276 5102 6328 5108
rect 5848 4380 6156 4389
rect 5848 4378 5854 4380
rect 5910 4378 5934 4380
rect 5990 4378 6014 4380
rect 6070 4378 6094 4380
rect 6150 4378 6156 4380
rect 5910 4326 5912 4378
rect 6092 4326 6094 4378
rect 5848 4324 5854 4326
rect 5910 4324 5934 4326
rect 5990 4324 6014 4326
rect 6070 4324 6094 4326
rect 6150 4324 6156 4326
rect 5848 4315 6156 4324
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5848 3292 6156 3301
rect 5848 3290 5854 3292
rect 5910 3290 5934 3292
rect 5990 3290 6014 3292
rect 6070 3290 6094 3292
rect 6150 3290 6156 3292
rect 5910 3238 5912 3290
rect 6092 3238 6094 3290
rect 5848 3236 5854 3238
rect 5910 3236 5934 3238
rect 5990 3236 6014 3238
rect 6070 3236 6094 3238
rect 6150 3236 6156 3238
rect 5848 3227 6156 3236
rect 6288 2990 6316 5102
rect 6656 3058 6684 6734
rect 6932 3534 6960 7754
rect 7208 7410 7236 8774
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7300 7750 7328 8434
rect 7576 7954 7604 8910
rect 8036 8294 8064 10678
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8128 8974 8156 10406
rect 8298 10364 8606 10373
rect 8298 10362 8304 10364
rect 8360 10362 8384 10364
rect 8440 10362 8464 10364
rect 8520 10362 8544 10364
rect 8600 10362 8606 10364
rect 8360 10310 8362 10362
rect 8542 10310 8544 10362
rect 8298 10308 8304 10310
rect 8360 10308 8384 10310
rect 8440 10308 8464 10310
rect 8520 10308 8544 10310
rect 8600 10308 8606 10310
rect 8298 10299 8606 10308
rect 8298 9276 8606 9285
rect 8298 9274 8304 9276
rect 8360 9274 8384 9276
rect 8440 9274 8464 9276
rect 8520 9274 8544 9276
rect 8600 9274 8606 9276
rect 8360 9222 8362 9274
rect 8542 9222 8544 9274
rect 8298 9220 8304 9222
rect 8360 9220 8384 9222
rect 8440 9220 8464 9222
rect 8520 9220 8544 9222
rect 8600 9220 8606 9222
rect 8298 9211 8606 9220
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 8036 7886 8064 8230
rect 8298 8188 8606 8197
rect 8298 8186 8304 8188
rect 8360 8186 8384 8188
rect 8440 8186 8464 8188
rect 8520 8186 8544 8188
rect 8600 8186 8606 8188
rect 8360 8134 8362 8186
rect 8542 8134 8544 8186
rect 8298 8132 8304 8134
rect 8360 8132 8384 8134
rect 8440 8132 8464 8134
rect 8520 8132 8544 8134
rect 8600 8132 8606 8134
rect 8298 8123 8606 8132
rect 8680 8090 8708 8366
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7300 7546 7328 7686
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 8220 7410 8248 7754
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8298 7100 8606 7109
rect 8298 7098 8304 7100
rect 8360 7098 8384 7100
rect 8440 7098 8464 7100
rect 8520 7098 8544 7100
rect 8600 7098 8606 7100
rect 8360 7046 8362 7098
rect 8542 7046 8544 7098
rect 8298 7044 8304 7046
rect 8360 7044 8384 7046
rect 8440 7044 8464 7046
rect 8520 7044 8544 7046
rect 8600 7044 8606 7046
rect 8298 7035 8606 7044
rect 8680 6798 8708 8026
rect 8772 6866 8800 19366
rect 8852 19304 8904 19310
rect 8852 19246 8904 19252
rect 8864 18426 8892 19246
rect 8852 18420 8904 18426
rect 8852 18362 8904 18368
rect 9048 18358 9076 19382
rect 9324 18630 9352 20810
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9600 20466 9628 20742
rect 9588 20460 9640 20466
rect 9588 20402 9640 20408
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9324 18426 9352 18566
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 9048 17610 9076 18294
rect 9036 17604 9088 17610
rect 9036 17546 9088 17552
rect 9324 16658 9352 18362
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 9232 15570 9260 15982
rect 9220 15564 9272 15570
rect 9220 15506 9272 15512
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 8956 12434 8984 12854
rect 9416 12434 9444 20334
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9692 18358 9720 19110
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 8956 12406 9076 12434
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 7748 6724 7800 6730
rect 7748 6666 7800 6672
rect 7024 6458 7052 6666
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 7024 5302 7052 5714
rect 7012 5296 7064 5302
rect 7012 5238 7064 5244
rect 7024 4622 7052 5238
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 7760 3738 7788 6666
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8298 6012 8606 6021
rect 8298 6010 8304 6012
rect 8360 6010 8384 6012
rect 8440 6010 8464 6012
rect 8520 6010 8544 6012
rect 8600 6010 8606 6012
rect 8360 5958 8362 6010
rect 8542 5958 8544 6010
rect 8298 5956 8304 5958
rect 8360 5956 8384 5958
rect 8440 5956 8464 5958
rect 8520 5956 8544 5958
rect 8600 5956 8606 5958
rect 8298 5947 8606 5956
rect 8680 5846 8708 6258
rect 8668 5840 8720 5846
rect 8668 5782 8720 5788
rect 8772 5710 8800 6598
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8668 5296 8720 5302
rect 8668 5238 8720 5244
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8220 4758 8248 4966
rect 8298 4924 8606 4933
rect 8298 4922 8304 4924
rect 8360 4922 8384 4924
rect 8440 4922 8464 4924
rect 8520 4922 8544 4924
rect 8600 4922 8606 4924
rect 8360 4870 8362 4922
rect 8542 4870 8544 4922
rect 8298 4868 8304 4870
rect 8360 4868 8384 4870
rect 8440 4868 8464 4870
rect 8520 4868 8544 4870
rect 8600 4868 8606 4870
rect 8298 4859 8606 4868
rect 8680 4826 8708 5238
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 7944 4146 7972 4558
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 8220 4078 8248 4694
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 7104 3392 7156 3398
rect 7760 3380 7788 3674
rect 8220 3602 8248 3878
rect 8298 3836 8606 3845
rect 8298 3834 8304 3836
rect 8360 3834 8384 3836
rect 8440 3834 8464 3836
rect 8520 3834 8544 3836
rect 8600 3834 8606 3836
rect 8360 3782 8362 3834
rect 8542 3782 8544 3834
rect 8298 3780 8304 3782
rect 8360 3780 8384 3782
rect 8440 3780 8464 3782
rect 8520 3780 8544 3782
rect 8600 3780 8606 3782
rect 8298 3771 8606 3780
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8680 3466 8708 4762
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 7104 3334 7156 3340
rect 7668 3352 7788 3380
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 4988 2508 5040 2514
rect 4988 2450 5040 2456
rect 4804 2372 4856 2378
rect 4804 2314 4856 2320
rect 5276 2310 5304 2926
rect 7116 2446 7144 3334
rect 7668 3126 7696 3352
rect 7656 3120 7708 3126
rect 7656 3062 7708 3068
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8298 2748 8606 2757
rect 8298 2746 8304 2748
rect 8360 2746 8384 2748
rect 8440 2746 8464 2748
rect 8520 2746 8544 2748
rect 8600 2746 8606 2748
rect 8360 2694 8362 2746
rect 8542 2694 8544 2746
rect 8298 2692 8304 2694
rect 8360 2692 8384 2694
rect 8440 2692 8464 2694
rect 8520 2692 8544 2694
rect 8600 2692 8606 2694
rect 8298 2683 8606 2692
rect 8680 2446 8708 2790
rect 8956 2514 8984 11290
rect 9048 8090 9076 12406
rect 9324 12406 9444 12434
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9232 10810 9260 11086
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9140 10266 9168 10542
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9324 9722 9352 12406
rect 9508 11354 9536 17070
rect 9600 16794 9628 17138
rect 9784 17134 9812 20878
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 9968 17882 9996 20470
rect 9956 17876 10008 17882
rect 9956 17818 10008 17824
rect 9968 17270 9996 17818
rect 10060 17338 10088 21490
rect 10508 20800 10560 20806
rect 10508 20742 10560 20748
rect 10324 19372 10376 19378
rect 10324 19314 10376 19320
rect 10336 18834 10364 19314
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 9956 17264 10008 17270
rect 9956 17206 10008 17212
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9784 16998 9812 17070
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9784 15586 9812 16934
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9876 16250 9904 16526
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9784 15558 9904 15586
rect 9680 15428 9732 15434
rect 9732 15388 9812 15416
rect 9680 15370 9732 15376
rect 9784 15162 9812 15388
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9600 13326 9628 13670
rect 9876 13326 9904 15558
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 9968 15094 9996 15302
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 10520 13530 10548 20742
rect 10747 20700 11055 20709
rect 10747 20698 10753 20700
rect 10809 20698 10833 20700
rect 10889 20698 10913 20700
rect 10969 20698 10993 20700
rect 11049 20698 11055 20700
rect 10809 20646 10811 20698
rect 10991 20646 10993 20698
rect 10747 20644 10753 20646
rect 10809 20644 10833 20646
rect 10889 20644 10913 20646
rect 10969 20644 10993 20646
rect 11049 20644 11055 20646
rect 10747 20635 11055 20644
rect 11624 20602 11652 21490
rect 12636 21146 12664 21490
rect 13197 21244 13505 21253
rect 13197 21242 13203 21244
rect 13259 21242 13283 21244
rect 13339 21242 13363 21244
rect 13419 21242 13443 21244
rect 13499 21242 13505 21244
rect 13259 21190 13261 21242
rect 13441 21190 13443 21242
rect 13197 21188 13203 21190
rect 13259 21188 13283 21190
rect 13339 21188 13363 21190
rect 13419 21188 13443 21190
rect 13499 21188 13505 21190
rect 13197 21179 13505 21188
rect 12624 21140 12676 21146
rect 12624 21082 12676 21088
rect 12532 20868 12584 20874
rect 12532 20810 12584 20816
rect 13084 20868 13136 20874
rect 13084 20810 13136 20816
rect 13820 20868 13872 20874
rect 13820 20810 13872 20816
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 11520 20392 11572 20398
rect 11520 20334 11572 20340
rect 11532 19854 11560 20334
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 10747 19612 11055 19621
rect 10747 19610 10753 19612
rect 10809 19610 10833 19612
rect 10889 19610 10913 19612
rect 10969 19610 10993 19612
rect 11049 19610 11055 19612
rect 10809 19558 10811 19610
rect 10991 19558 10993 19610
rect 10747 19556 10753 19558
rect 10809 19556 10833 19558
rect 10889 19556 10913 19558
rect 10969 19556 10993 19558
rect 11049 19556 11055 19558
rect 10747 19547 11055 19556
rect 11532 19378 11560 19790
rect 12440 19780 12492 19786
rect 12440 19722 12492 19728
rect 12452 19514 12480 19722
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11796 19304 11848 19310
rect 11796 19246 11848 19252
rect 11808 18970 11836 19246
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 10600 18692 10652 18698
rect 10600 18634 10652 18640
rect 10612 18426 10640 18634
rect 10747 18524 11055 18533
rect 10747 18522 10753 18524
rect 10809 18522 10833 18524
rect 10889 18522 10913 18524
rect 10969 18522 10993 18524
rect 11049 18522 11055 18524
rect 10809 18470 10811 18522
rect 10991 18470 10993 18522
rect 10747 18468 10753 18470
rect 10809 18468 10833 18470
rect 10889 18468 10913 18470
rect 10969 18468 10993 18470
rect 11049 18468 11055 18470
rect 10747 18459 11055 18468
rect 10600 18420 10652 18426
rect 10600 18362 10652 18368
rect 12544 17610 12572 20810
rect 12808 20528 12860 20534
rect 12808 20470 12860 20476
rect 12820 19718 12848 20470
rect 13096 20398 13124 20810
rect 13084 20392 13136 20398
rect 13084 20334 13136 20340
rect 13197 20156 13505 20165
rect 13197 20154 13203 20156
rect 13259 20154 13283 20156
rect 13339 20154 13363 20156
rect 13419 20154 13443 20156
rect 13499 20154 13505 20156
rect 13259 20102 13261 20154
rect 13441 20102 13443 20154
rect 13197 20100 13203 20102
rect 13259 20100 13283 20102
rect 13339 20100 13363 20102
rect 13419 20100 13443 20102
rect 13499 20100 13505 20102
rect 13197 20091 13505 20100
rect 13832 19718 13860 20810
rect 13912 20392 13964 20398
rect 13912 20334 13964 20340
rect 13924 20058 13952 20334
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 12820 19446 12848 19654
rect 12808 19440 12860 19446
rect 12808 19382 12860 19388
rect 12820 18630 12848 19382
rect 13197 19068 13505 19077
rect 13197 19066 13203 19068
rect 13259 19066 13283 19068
rect 13339 19066 13363 19068
rect 13419 19066 13443 19068
rect 13499 19066 13505 19068
rect 13259 19014 13261 19066
rect 13441 19014 13443 19066
rect 13197 19012 13203 19014
rect 13259 19012 13283 19014
rect 13339 19012 13363 19014
rect 13419 19012 13443 19014
rect 13499 19012 13505 19014
rect 13197 19003 13505 19012
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12532 17604 12584 17610
rect 12532 17546 12584 17552
rect 11244 17536 11296 17542
rect 11244 17478 11296 17484
rect 10747 17436 11055 17445
rect 10747 17434 10753 17436
rect 10809 17434 10833 17436
rect 10889 17434 10913 17436
rect 10969 17434 10993 17436
rect 11049 17434 11055 17436
rect 10809 17382 10811 17434
rect 10991 17382 10993 17434
rect 10747 17380 10753 17382
rect 10809 17380 10833 17382
rect 10889 17380 10913 17382
rect 10969 17380 10993 17382
rect 11049 17380 11055 17382
rect 10747 17371 11055 17380
rect 11256 17338 11284 17478
rect 11244 17332 11296 17338
rect 11244 17274 11296 17280
rect 10747 16348 11055 16357
rect 10747 16346 10753 16348
rect 10809 16346 10833 16348
rect 10889 16346 10913 16348
rect 10969 16346 10993 16348
rect 11049 16346 11055 16348
rect 10809 16294 10811 16346
rect 10991 16294 10993 16346
rect 10747 16292 10753 16294
rect 10809 16292 10833 16294
rect 10889 16292 10913 16294
rect 10969 16292 10993 16294
rect 11049 16292 11055 16294
rect 10747 16283 11055 16292
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11256 15706 11284 16050
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 10747 15260 11055 15269
rect 10747 15258 10753 15260
rect 10809 15258 10833 15260
rect 10889 15258 10913 15260
rect 10969 15258 10993 15260
rect 11049 15258 11055 15260
rect 10809 15206 10811 15258
rect 10991 15206 10993 15258
rect 10747 15204 10753 15206
rect 10809 15204 10833 15206
rect 10889 15204 10913 15206
rect 10969 15204 10993 15206
rect 11049 15204 11055 15206
rect 10747 15195 11055 15204
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11164 14822 11192 14962
rect 11624 14958 11652 15438
rect 12440 15428 12492 15434
rect 12440 15370 12492 15376
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 10747 14172 11055 14181
rect 10747 14170 10753 14172
rect 10809 14170 10833 14172
rect 10889 14170 10913 14172
rect 10969 14170 10993 14172
rect 11049 14170 11055 14172
rect 10809 14118 10811 14170
rect 10991 14118 10993 14170
rect 10747 14116 10753 14118
rect 10809 14116 10833 14118
rect 10889 14116 10913 14118
rect 10969 14116 10993 14118
rect 11049 14116 11055 14118
rect 10747 14107 11055 14116
rect 11164 13802 11192 14758
rect 11152 13796 11204 13802
rect 11152 13738 11204 13744
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10324 13184 10376 13190
rect 10324 13126 10376 13132
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9876 12434 9904 12582
rect 9876 12406 9996 12434
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9140 7410 9168 7686
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9324 3058 9352 9658
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9508 7478 9536 8230
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9508 6322 9536 7414
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9600 5234 9628 6054
rect 9692 5658 9720 10678
rect 9784 10606 9812 11086
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9876 10266 9904 11086
rect 9968 11082 9996 12406
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 10060 10266 10088 10406
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10244 10130 10272 12786
rect 10336 12782 10364 13126
rect 10428 12850 10456 13262
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 10520 12434 10548 13466
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 10600 13252 10652 13258
rect 10600 13194 10652 13200
rect 10612 12782 10640 13194
rect 10747 13084 11055 13093
rect 10747 13082 10753 13084
rect 10809 13082 10833 13084
rect 10889 13082 10913 13084
rect 10969 13082 10993 13084
rect 11049 13082 11055 13084
rect 10809 13030 10811 13082
rect 10991 13030 10993 13082
rect 10747 13028 10753 13030
rect 10809 13028 10833 13030
rect 10889 13028 10913 13030
rect 10969 13028 10993 13030
rect 11049 13028 11055 13030
rect 10747 13019 11055 13028
rect 11992 12986 12020 13262
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 12176 12850 12204 13330
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 11060 12708 11112 12714
rect 11060 12650 11112 12656
rect 11072 12442 11100 12650
rect 11060 12436 11112 12442
rect 10520 12406 10640 12434
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10520 10062 10548 10406
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10508 8288 10560 8294
rect 10508 8230 10560 8236
rect 10520 7818 10548 8230
rect 10416 7812 10468 7818
rect 10416 7754 10468 7760
rect 10508 7812 10560 7818
rect 10508 7754 10560 7760
rect 10428 7546 10456 7754
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10520 7410 10548 7754
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10508 7268 10560 7274
rect 10508 7210 10560 7216
rect 10520 6662 10548 7210
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10520 5778 10548 6598
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 9692 5642 9812 5658
rect 9692 5636 9824 5642
rect 9692 5630 9772 5636
rect 9772 5578 9824 5584
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9784 3534 9812 5578
rect 10508 5092 10560 5098
rect 10508 5034 10560 5040
rect 10520 4690 10548 5034
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 10612 3602 10640 12406
rect 11060 12378 11112 12384
rect 12452 12170 12480 15370
rect 12544 13802 12572 17546
rect 12820 16794 12848 18566
rect 13197 17980 13505 17989
rect 13197 17978 13203 17980
rect 13259 17978 13283 17980
rect 13339 17978 13363 17980
rect 13419 17978 13443 17980
rect 13499 17978 13505 17980
rect 13259 17926 13261 17978
rect 13441 17926 13443 17978
rect 13197 17924 13203 17926
rect 13259 17924 13283 17926
rect 13339 17924 13363 17926
rect 13419 17924 13443 17926
rect 13499 17924 13505 17926
rect 13197 17915 13505 17924
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13556 17270 13584 17614
rect 13544 17264 13596 17270
rect 13544 17206 13596 17212
rect 13740 17134 13768 17682
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14108 17202 14136 17614
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13197 16892 13505 16901
rect 13197 16890 13203 16892
rect 13259 16890 13283 16892
rect 13339 16890 13363 16892
rect 13419 16890 13443 16892
rect 13499 16890 13505 16892
rect 13259 16838 13261 16890
rect 13441 16838 13443 16890
rect 13197 16836 13203 16838
rect 13259 16836 13283 16838
rect 13339 16836 13363 16838
rect 13419 16836 13443 16838
rect 13499 16836 13505 16838
rect 13197 16827 13505 16836
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 13197 15804 13505 15813
rect 13197 15802 13203 15804
rect 13259 15802 13283 15804
rect 13339 15802 13363 15804
rect 13419 15802 13443 15804
rect 13499 15802 13505 15804
rect 13259 15750 13261 15802
rect 13441 15750 13443 15802
rect 13197 15748 13203 15750
rect 13259 15748 13283 15750
rect 13339 15748 13363 15750
rect 13419 15748 13443 15750
rect 13499 15748 13505 15750
rect 13197 15739 13505 15748
rect 14200 15706 14228 21490
rect 14372 20868 14424 20874
rect 14372 20810 14424 20816
rect 14384 20602 14412 20810
rect 14372 20596 14424 20602
rect 14372 20538 14424 20544
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14384 17338 14412 18226
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 14924 17196 14976 17202
rect 14924 17138 14976 17144
rect 14936 15910 14964 17138
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14372 15632 14424 15638
rect 14372 15574 14424 15580
rect 13268 15428 13320 15434
rect 13268 15370 13320 15376
rect 13280 15094 13308 15370
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 14004 15088 14056 15094
rect 14004 15030 14056 15036
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13197 14716 13505 14725
rect 13197 14714 13203 14716
rect 13259 14714 13283 14716
rect 13339 14714 13363 14716
rect 13419 14714 13443 14716
rect 13499 14714 13505 14716
rect 13259 14662 13261 14714
rect 13441 14662 13443 14714
rect 13197 14660 13203 14662
rect 13259 14660 13283 14662
rect 13339 14660 13363 14662
rect 13419 14660 13443 14662
rect 13499 14660 13505 14662
rect 13197 14651 13505 14660
rect 13924 14482 13952 14894
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 12544 13462 12572 13738
rect 13096 13530 13124 13874
rect 13197 13628 13505 13637
rect 13197 13626 13203 13628
rect 13259 13626 13283 13628
rect 13339 13626 13363 13628
rect 13419 13626 13443 13628
rect 13499 13626 13505 13628
rect 13259 13574 13261 13626
rect 13441 13574 13443 13626
rect 13197 13572 13203 13574
rect 13259 13572 13283 13574
rect 13339 13572 13363 13574
rect 13419 13572 13443 13574
rect 13499 13572 13505 13574
rect 13197 13563 13505 13572
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 13924 13394 13952 14418
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12544 12986 12572 13262
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 13197 12540 13505 12549
rect 13197 12538 13203 12540
rect 13259 12538 13283 12540
rect 13339 12538 13363 12540
rect 13419 12538 13443 12540
rect 13499 12538 13505 12540
rect 13259 12486 13261 12538
rect 13441 12486 13443 12538
rect 13197 12484 13203 12486
rect 13259 12484 13283 12486
rect 13339 12484 13363 12486
rect 13419 12484 13443 12486
rect 13499 12484 13505 12486
rect 13197 12475 13505 12484
rect 13924 12306 13952 13330
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 10747 11996 11055 12005
rect 10747 11994 10753 11996
rect 10809 11994 10833 11996
rect 10889 11994 10913 11996
rect 10969 11994 10993 11996
rect 11049 11994 11055 11996
rect 10809 11942 10811 11994
rect 10991 11942 10993 11994
rect 10747 11940 10753 11942
rect 10809 11940 10833 11942
rect 10889 11940 10913 11942
rect 10969 11940 10993 11942
rect 11049 11940 11055 11942
rect 10747 11931 11055 11940
rect 12452 11898 12480 12106
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11716 11354 11744 11630
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 10747 10908 11055 10917
rect 10747 10906 10753 10908
rect 10809 10906 10833 10908
rect 10889 10906 10913 10908
rect 10969 10906 10993 10908
rect 11049 10906 11055 10908
rect 10809 10854 10811 10906
rect 10991 10854 10993 10906
rect 10747 10852 10753 10854
rect 10809 10852 10833 10854
rect 10889 10852 10913 10854
rect 10969 10852 10993 10854
rect 11049 10852 11055 10854
rect 10747 10843 11055 10852
rect 11164 10810 11192 11086
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10980 10062 11008 10542
rect 11256 10130 11284 10746
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10747 9820 11055 9829
rect 10747 9818 10753 9820
rect 10809 9818 10833 9820
rect 10889 9818 10913 9820
rect 10969 9818 10993 9820
rect 11049 9818 11055 9820
rect 10809 9766 10811 9818
rect 10991 9766 10993 9818
rect 10747 9764 10753 9766
rect 10809 9764 10833 9766
rect 10889 9764 10913 9766
rect 10969 9764 10993 9766
rect 11049 9764 11055 9766
rect 10747 9755 11055 9764
rect 10747 8732 11055 8741
rect 10747 8730 10753 8732
rect 10809 8730 10833 8732
rect 10889 8730 10913 8732
rect 10969 8730 10993 8732
rect 11049 8730 11055 8732
rect 10809 8678 10811 8730
rect 10991 8678 10993 8730
rect 10747 8676 10753 8678
rect 10809 8676 10833 8678
rect 10889 8676 10913 8678
rect 10969 8676 10993 8678
rect 11049 8676 11055 8678
rect 10747 8667 11055 8676
rect 10747 7644 11055 7653
rect 10747 7642 10753 7644
rect 10809 7642 10833 7644
rect 10889 7642 10913 7644
rect 10969 7642 10993 7644
rect 11049 7642 11055 7644
rect 10809 7590 10811 7642
rect 10991 7590 10993 7642
rect 10747 7588 10753 7590
rect 10809 7588 10833 7590
rect 10889 7588 10913 7590
rect 10969 7588 10993 7590
rect 11049 7588 11055 7590
rect 10747 7579 11055 7588
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10980 6798 11008 7142
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 11256 6610 11284 10066
rect 11440 10062 11468 11154
rect 11808 10810 11836 11630
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11532 9926 11560 10610
rect 11900 10470 11928 11698
rect 13197 11452 13505 11461
rect 13197 11450 13203 11452
rect 13259 11450 13283 11452
rect 13339 11450 13363 11452
rect 13419 11450 13443 11452
rect 13499 11450 13505 11452
rect 13259 11398 13261 11450
rect 13441 11398 13443 11450
rect 13197 11396 13203 11398
rect 13259 11396 13283 11398
rect 13339 11396 13363 11398
rect 13419 11396 13443 11398
rect 13499 11396 13505 11398
rect 13197 11387 13505 11396
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12176 9994 12204 10406
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 12360 9586 12388 11154
rect 13197 10364 13505 10373
rect 13197 10362 13203 10364
rect 13259 10362 13283 10364
rect 13339 10362 13363 10364
rect 13419 10362 13443 10364
rect 13499 10362 13505 10364
rect 13259 10310 13261 10362
rect 13441 10310 13443 10362
rect 13197 10308 13203 10310
rect 13259 10308 13283 10310
rect 13339 10308 13363 10310
rect 13419 10308 13443 10310
rect 13499 10308 13505 10310
rect 13197 10299 13505 10308
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 13096 9722 13124 10066
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13188 9586 13216 10134
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13556 9722 13584 9998
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13197 9276 13505 9285
rect 13197 9274 13203 9276
rect 13259 9274 13283 9276
rect 13339 9274 13363 9276
rect 13419 9274 13443 9276
rect 13499 9274 13505 9276
rect 13259 9222 13261 9274
rect 13441 9222 13443 9274
rect 13197 9220 13203 9222
rect 13259 9220 13283 9222
rect 13339 9220 13363 9222
rect 13419 9220 13443 9222
rect 13499 9220 13505 9222
rect 13197 9211 13505 9220
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11808 7478 11836 8230
rect 11900 8090 11928 8434
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11992 7954 12020 8230
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 12452 7546 12480 8434
rect 12544 7750 12572 8434
rect 13197 8188 13505 8197
rect 13197 8186 13203 8188
rect 13259 8186 13283 8188
rect 13339 8186 13363 8188
rect 13419 8186 13443 8188
rect 13499 8186 13505 8188
rect 13259 8134 13261 8186
rect 13441 8134 13443 8186
rect 13197 8132 13203 8134
rect 13259 8132 13283 8134
rect 13339 8132 13363 8134
rect 13419 8132 13443 8134
rect 13499 8132 13505 8134
rect 13197 8123 13505 8132
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 11796 7472 11848 7478
rect 11796 7414 11848 7420
rect 12544 7342 12572 7686
rect 12728 7546 12756 7754
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11256 6582 11376 6610
rect 10747 6556 11055 6565
rect 10747 6554 10753 6556
rect 10809 6554 10833 6556
rect 10889 6554 10913 6556
rect 10969 6554 10993 6556
rect 11049 6554 11055 6556
rect 10809 6502 10811 6554
rect 10991 6502 10993 6554
rect 10747 6500 10753 6502
rect 10809 6500 10833 6502
rect 10889 6500 10913 6502
rect 10969 6500 10993 6502
rect 11049 6500 11055 6502
rect 10747 6491 11055 6500
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11256 5710 11284 6394
rect 11348 5778 11376 6582
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 10747 5468 11055 5477
rect 10747 5466 10753 5468
rect 10809 5466 10833 5468
rect 10889 5466 10913 5468
rect 10969 5466 10993 5468
rect 11049 5466 11055 5468
rect 10809 5414 10811 5466
rect 10991 5414 10993 5466
rect 10747 5412 10753 5414
rect 10809 5412 10833 5414
rect 10889 5412 10913 5414
rect 10969 5412 10993 5414
rect 11049 5412 11055 5414
rect 10747 5403 11055 5412
rect 11348 4690 11376 5714
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 10747 4380 11055 4389
rect 10747 4378 10753 4380
rect 10809 4378 10833 4380
rect 10889 4378 10913 4380
rect 10969 4378 10993 4380
rect 11049 4378 11055 4380
rect 10809 4326 10811 4378
rect 10991 4326 10993 4378
rect 10747 4324 10753 4326
rect 10809 4324 10833 4326
rect 10889 4324 10913 4326
rect 10969 4324 10993 4326
rect 11049 4324 11055 4326
rect 10747 4315 11055 4324
rect 11348 3602 11376 4626
rect 11900 4010 11928 7142
rect 13197 7100 13505 7109
rect 13197 7098 13203 7100
rect 13259 7098 13283 7100
rect 13339 7098 13363 7100
rect 13419 7098 13443 7100
rect 13499 7098 13505 7100
rect 13259 7046 13261 7098
rect 13441 7046 13443 7098
rect 13197 7044 13203 7046
rect 13259 7044 13283 7046
rect 13339 7044 13363 7046
rect 13419 7044 13443 7046
rect 13499 7044 13505 7046
rect 13197 7035 13505 7044
rect 13648 6914 13676 12038
rect 13924 11914 13952 12242
rect 13832 11898 13952 11914
rect 13820 11892 13952 11898
rect 13872 11886 13952 11892
rect 13820 11834 13872 11840
rect 14016 11830 14044 15030
rect 14292 14346 14320 15302
rect 14280 14340 14332 14346
rect 14280 14282 14332 14288
rect 14384 13394 14412 15574
rect 14936 15570 14964 15846
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 14556 15428 14608 15434
rect 14556 15370 14608 15376
rect 14568 13938 14596 15370
rect 15028 15162 15056 21490
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 15212 19922 15240 20742
rect 15396 19938 15424 20946
rect 15646 20700 15954 20709
rect 15646 20698 15652 20700
rect 15708 20698 15732 20700
rect 15788 20698 15812 20700
rect 15868 20698 15892 20700
rect 15948 20698 15954 20700
rect 15708 20646 15710 20698
rect 15890 20646 15892 20698
rect 15646 20644 15652 20646
rect 15708 20644 15732 20646
rect 15788 20644 15812 20646
rect 15868 20644 15892 20646
rect 15948 20644 15954 20646
rect 15646 20635 15954 20644
rect 16488 20256 16540 20262
rect 16488 20198 16540 20204
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 15304 19910 15424 19938
rect 15304 19854 15332 19910
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15580 18086 15608 19790
rect 15646 19612 15954 19621
rect 15646 19610 15652 19612
rect 15708 19610 15732 19612
rect 15788 19610 15812 19612
rect 15868 19610 15892 19612
rect 15948 19610 15954 19612
rect 15708 19558 15710 19610
rect 15890 19558 15892 19610
rect 15646 19556 15652 19558
rect 15708 19556 15732 19558
rect 15788 19556 15812 19558
rect 15868 19556 15892 19558
rect 15948 19556 15954 19558
rect 15646 19547 15954 19556
rect 16028 18760 16080 18766
rect 16028 18702 16080 18708
rect 15646 18524 15954 18533
rect 15646 18522 15652 18524
rect 15708 18522 15732 18524
rect 15788 18522 15812 18524
rect 15868 18522 15892 18524
rect 15948 18522 15954 18524
rect 15708 18470 15710 18522
rect 15890 18470 15892 18522
rect 15646 18468 15652 18470
rect 15708 18468 15732 18470
rect 15788 18468 15812 18470
rect 15868 18468 15892 18470
rect 15948 18468 15954 18470
rect 15646 18459 15954 18468
rect 16040 18426 16068 18702
rect 16028 18420 16080 18426
rect 16028 18362 16080 18368
rect 15660 18352 15712 18358
rect 15660 18294 15712 18300
rect 15672 18154 15700 18294
rect 15660 18148 15712 18154
rect 15660 18090 15712 18096
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 14384 12714 14412 13330
rect 14568 12986 14596 13874
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 14372 12708 14424 12714
rect 14372 12650 14424 12656
rect 14648 12708 14700 12714
rect 14648 12650 14700 12656
rect 14660 12306 14688 12650
rect 14648 12300 14700 12306
rect 14648 12242 14700 12248
rect 14660 12170 14688 12242
rect 15120 12170 15148 12922
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 15108 12164 15160 12170
rect 15108 12106 15160 12112
rect 14004 11824 14056 11830
rect 14004 11766 14056 11772
rect 14016 11354 14044 11766
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14108 10810 14136 11086
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14476 10266 14504 10610
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13740 9450 13768 9998
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14292 7954 14320 8230
rect 14280 7948 14332 7954
rect 14280 7890 14332 7896
rect 14740 7812 14792 7818
rect 14740 7754 14792 7760
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 13924 7342 13952 7686
rect 14108 7546 14136 7686
rect 14752 7546 14780 7754
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 13556 6886 13676 6914
rect 13197 6012 13505 6021
rect 13197 6010 13203 6012
rect 13259 6010 13283 6012
rect 13339 6010 13363 6012
rect 13419 6010 13443 6012
rect 13499 6010 13505 6012
rect 13259 5958 13261 6010
rect 13441 5958 13443 6010
rect 13197 5956 13203 5958
rect 13259 5956 13283 5958
rect 13339 5956 13363 5958
rect 13419 5956 13443 5958
rect 13499 5956 13505 5958
rect 13197 5947 13505 5956
rect 12164 5636 12216 5642
rect 12164 5578 12216 5584
rect 12176 4554 12204 5578
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12268 4826 12296 5170
rect 13197 4924 13505 4933
rect 13197 4922 13203 4924
rect 13259 4922 13283 4924
rect 13339 4922 13363 4924
rect 13419 4922 13443 4924
rect 13499 4922 13505 4924
rect 13259 4870 13261 4922
rect 13441 4870 13443 4922
rect 13197 4868 13203 4870
rect 13259 4868 13283 4870
rect 13339 4868 13363 4870
rect 13419 4868 13443 4870
rect 13499 4868 13505 4870
rect 13197 4859 13505 4868
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 12176 4026 12204 4490
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 12084 3998 12204 4026
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9508 2514 9536 2926
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 5736 800 5764 2246
rect 5848 2204 6156 2213
rect 5848 2202 5854 2204
rect 5910 2202 5934 2204
rect 5990 2202 6014 2204
rect 6070 2202 6094 2204
rect 6150 2202 6156 2204
rect 5910 2150 5912 2202
rect 6092 2150 6094 2202
rect 5848 2148 5854 2150
rect 5910 2148 5934 2150
rect 5990 2148 6014 2150
rect 6070 2148 6094 2150
rect 6150 2148 6156 2150
rect 5848 2139 6156 2148
rect 7024 800 7052 2246
rect 8312 800 8340 2246
rect 9600 800 9628 3334
rect 10244 3126 10272 3334
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 10336 2650 10364 3470
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10520 2378 10548 3470
rect 10747 3292 11055 3301
rect 10747 3290 10753 3292
rect 10809 3290 10833 3292
rect 10889 3290 10913 3292
rect 10969 3290 10993 3292
rect 11049 3290 11055 3292
rect 10809 3238 10811 3290
rect 10991 3238 10993 3290
rect 10747 3236 10753 3238
rect 10809 3236 10833 3238
rect 10889 3236 10913 3238
rect 10969 3236 10993 3238
rect 11049 3236 11055 3238
rect 10747 3227 11055 3236
rect 11348 2922 11376 3538
rect 11900 2990 11928 3946
rect 12084 3466 12112 3998
rect 13197 3836 13505 3845
rect 13197 3834 13203 3836
rect 13259 3834 13283 3836
rect 13339 3834 13363 3836
rect 13419 3834 13443 3836
rect 13499 3834 13505 3836
rect 13259 3782 13261 3834
rect 13441 3782 13443 3834
rect 13197 3780 13203 3782
rect 13259 3780 13283 3782
rect 13339 3780 13363 3782
rect 13419 3780 13443 3782
rect 13499 3780 13505 3782
rect 13197 3771 13505 3780
rect 12072 3460 12124 3466
rect 12072 3402 12124 3408
rect 12084 3126 12112 3402
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 11336 2916 11388 2922
rect 11336 2858 11388 2864
rect 11244 2848 11296 2854
rect 11244 2790 11296 2796
rect 10600 2576 10652 2582
rect 10600 2518 10652 2524
rect 10508 2372 10560 2378
rect 10508 2314 10560 2320
rect 570 0 626 800
rect 1858 0 1914 800
rect 3146 0 3202 800
rect 4434 0 4490 800
rect 5722 0 5778 800
rect 7010 0 7066 800
rect 8298 0 8354 800
rect 9586 0 9642 800
rect 10612 762 10640 2518
rect 11256 2446 11284 2790
rect 12544 2446 12572 3334
rect 13197 2748 13505 2757
rect 13197 2746 13203 2748
rect 13259 2746 13283 2748
rect 13339 2746 13363 2748
rect 13419 2746 13443 2748
rect 13499 2746 13505 2748
rect 13259 2694 13261 2746
rect 13441 2694 13443 2746
rect 13197 2692 13203 2694
rect 13259 2692 13283 2694
rect 13339 2692 13363 2694
rect 13419 2692 13443 2694
rect 13499 2692 13505 2694
rect 13197 2683 13505 2692
rect 13556 2446 13584 6886
rect 13924 6798 13952 7278
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 14464 5840 14516 5846
rect 14464 5782 14516 5788
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13832 4622 13860 5510
rect 14096 5092 14148 5098
rect 14096 5034 14148 5040
rect 14108 4826 14136 5034
rect 14384 5030 14412 5714
rect 14476 5370 14504 5782
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14384 4690 14412 4966
rect 14372 4684 14424 4690
rect 14372 4626 14424 4632
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 15028 2446 15056 11494
rect 15108 4752 15160 4758
rect 15108 4694 15160 4700
rect 15120 3194 15148 4694
rect 15304 3602 15332 18022
rect 15672 17882 15700 18090
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 16500 17678 16528 20198
rect 16684 19786 16712 20198
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 16684 18850 16712 19722
rect 16592 18822 16712 18850
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 15646 17436 15954 17445
rect 15646 17434 15652 17436
rect 15708 17434 15732 17436
rect 15788 17434 15812 17436
rect 15868 17434 15892 17436
rect 15948 17434 15954 17436
rect 15708 17382 15710 17434
rect 15890 17382 15892 17434
rect 15646 17380 15652 17382
rect 15708 17380 15732 17382
rect 15788 17380 15812 17382
rect 15868 17380 15892 17382
rect 15948 17380 15954 17382
rect 15646 17371 15954 17380
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15488 16810 15516 17138
rect 15660 16992 15712 16998
rect 15660 16934 15712 16940
rect 15396 16782 15516 16810
rect 15396 16658 15424 16782
rect 15672 16658 15700 16934
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15396 15706 15424 16594
rect 16592 16454 16620 18822
rect 16776 16574 16804 21490
rect 17040 20936 17092 20942
rect 17040 20878 17092 20884
rect 17052 17338 17080 20878
rect 17512 20058 17540 21490
rect 18096 21244 18404 21253
rect 18096 21242 18102 21244
rect 18158 21242 18182 21244
rect 18238 21242 18262 21244
rect 18318 21242 18342 21244
rect 18398 21242 18404 21244
rect 18158 21190 18160 21242
rect 18340 21190 18342 21242
rect 18096 21188 18102 21190
rect 18158 21188 18182 21190
rect 18238 21188 18262 21190
rect 18318 21188 18342 21190
rect 18398 21188 18404 21190
rect 18096 21179 18404 21188
rect 19352 21146 19380 21490
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19628 20942 19656 21519
rect 19708 21490 19760 21496
rect 19616 20936 19668 20942
rect 19616 20878 19668 20884
rect 18972 20868 19024 20874
rect 18972 20810 19024 20816
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 18340 20346 18368 20402
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 17972 19378 18000 20334
rect 18340 20318 18460 20346
rect 18096 20156 18404 20165
rect 18096 20154 18102 20156
rect 18158 20154 18182 20156
rect 18238 20154 18262 20156
rect 18318 20154 18342 20156
rect 18398 20154 18404 20156
rect 18158 20102 18160 20154
rect 18340 20102 18342 20154
rect 18096 20100 18102 20102
rect 18158 20100 18182 20102
rect 18238 20100 18262 20102
rect 18318 20100 18342 20102
rect 18398 20100 18404 20102
rect 18096 20091 18404 20100
rect 18432 19854 18460 20318
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 18248 19446 18276 19654
rect 18236 19440 18288 19446
rect 18236 19382 18288 19388
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 17592 18760 17644 18766
rect 17592 18702 17644 18708
rect 17604 17746 17632 18702
rect 17972 18306 18000 19314
rect 18096 19068 18404 19077
rect 18096 19066 18102 19068
rect 18158 19066 18182 19068
rect 18238 19066 18262 19068
rect 18318 19066 18342 19068
rect 18398 19066 18404 19068
rect 18158 19014 18160 19066
rect 18340 19014 18342 19066
rect 18096 19012 18102 19014
rect 18158 19012 18182 19014
rect 18238 19012 18262 19014
rect 18318 19012 18342 19014
rect 18398 19012 18404 19014
rect 18096 19003 18404 19012
rect 18432 18358 18460 19790
rect 18788 19440 18840 19446
rect 18788 19382 18840 19388
rect 18800 18766 18828 19382
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18800 18358 18828 18702
rect 17880 18290 18000 18306
rect 18420 18352 18472 18358
rect 18420 18294 18472 18300
rect 18788 18352 18840 18358
rect 18788 18294 18840 18300
rect 17868 18284 18000 18290
rect 17920 18278 18000 18284
rect 17868 18226 17920 18232
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 17224 17332 17276 17338
rect 17224 17274 17276 17280
rect 17132 17060 17184 17066
rect 17132 17002 17184 17008
rect 17144 16794 17172 17002
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 17144 16590 17172 16730
rect 16684 16546 16804 16574
rect 17132 16584 17184 16590
rect 16580 16448 16632 16454
rect 16580 16390 16632 16396
rect 15646 16348 15954 16357
rect 15646 16346 15652 16348
rect 15708 16346 15732 16348
rect 15788 16346 15812 16348
rect 15868 16346 15892 16348
rect 15948 16346 15954 16348
rect 15708 16294 15710 16346
rect 15890 16294 15892 16346
rect 15646 16292 15652 16294
rect 15708 16292 15732 16294
rect 15788 16292 15812 16294
rect 15868 16292 15892 16294
rect 15948 16292 15954 16294
rect 15646 16283 15954 16292
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 16684 15450 16712 16546
rect 17236 16574 17264 17274
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17512 16794 17540 17138
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17604 16574 17632 17682
rect 17972 17542 18000 18278
rect 18096 17980 18404 17989
rect 18096 17978 18102 17980
rect 18158 17978 18182 17980
rect 18238 17978 18262 17980
rect 18318 17978 18342 17980
rect 18398 17978 18404 17980
rect 18158 17926 18160 17978
rect 18340 17926 18342 17978
rect 18096 17924 18102 17926
rect 18158 17924 18182 17926
rect 18238 17924 18262 17926
rect 18318 17924 18342 17926
rect 18398 17924 18404 17926
rect 18096 17915 18404 17924
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 17684 17264 17736 17270
rect 17684 17206 17736 17212
rect 17236 16546 17356 16574
rect 17132 16526 17184 16532
rect 17132 15564 17184 15570
rect 17132 15506 17184 15512
rect 16592 15422 16712 15450
rect 15646 15260 15954 15269
rect 15646 15258 15652 15260
rect 15708 15258 15732 15260
rect 15788 15258 15812 15260
rect 15868 15258 15892 15260
rect 15948 15258 15954 15260
rect 15708 15206 15710 15258
rect 15890 15206 15892 15258
rect 15646 15204 15652 15206
rect 15708 15204 15732 15206
rect 15788 15204 15812 15206
rect 15868 15204 15892 15206
rect 15948 15204 15954 15206
rect 15646 15195 15954 15204
rect 16592 14618 16620 15422
rect 17040 14884 17092 14890
rect 17040 14826 17092 14832
rect 17052 14618 17080 14826
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 17144 14414 17172 15506
rect 17224 14544 17276 14550
rect 17224 14486 17276 14492
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 15396 13870 15424 14282
rect 15646 14172 15954 14181
rect 15646 14170 15652 14172
rect 15708 14170 15732 14172
rect 15788 14170 15812 14172
rect 15868 14170 15892 14172
rect 15948 14170 15954 14172
rect 15708 14118 15710 14170
rect 15890 14118 15892 14170
rect 15646 14116 15652 14118
rect 15708 14116 15732 14118
rect 15788 14116 15812 14118
rect 15868 14116 15892 14118
rect 15948 14116 15954 14118
rect 15646 14107 15954 14116
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15396 13258 15424 13806
rect 15384 13252 15436 13258
rect 15384 13194 15436 13200
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 15646 13084 15954 13093
rect 15646 13082 15652 13084
rect 15708 13082 15732 13084
rect 15788 13082 15812 13084
rect 15868 13082 15892 13084
rect 15948 13082 15954 13084
rect 15708 13030 15710 13082
rect 15890 13030 15892 13082
rect 15646 13028 15652 13030
rect 15708 13028 15732 13030
rect 15788 13028 15812 13030
rect 15868 13028 15892 13030
rect 15948 13028 15954 13030
rect 15646 13019 15954 13028
rect 15646 11996 15954 12005
rect 15646 11994 15652 11996
rect 15708 11994 15732 11996
rect 15788 11994 15812 11996
rect 15868 11994 15892 11996
rect 15948 11994 15954 11996
rect 15708 11942 15710 11994
rect 15890 11942 15892 11994
rect 15646 11940 15652 11942
rect 15708 11940 15732 11942
rect 15788 11940 15812 11942
rect 15868 11940 15892 11942
rect 15948 11940 15954 11942
rect 15646 11931 15954 11940
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15672 11218 15700 11630
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15384 11008 15436 11014
rect 15384 10950 15436 10956
rect 15396 9926 15424 10950
rect 15646 10908 15954 10917
rect 15646 10906 15652 10908
rect 15708 10906 15732 10908
rect 15788 10906 15812 10908
rect 15868 10906 15892 10908
rect 15948 10906 15954 10908
rect 15708 10854 15710 10906
rect 15890 10854 15892 10906
rect 15646 10852 15652 10854
rect 15708 10852 15732 10854
rect 15788 10852 15812 10854
rect 15868 10852 15892 10854
rect 15948 10852 15954 10854
rect 15646 10843 15954 10852
rect 16040 10010 16068 13126
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16408 12170 16436 12310
rect 16396 12164 16448 12170
rect 16396 12106 16448 12112
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 16040 9982 16160 10010
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15396 6118 15424 9862
rect 15646 9820 15954 9829
rect 15646 9818 15652 9820
rect 15708 9818 15732 9820
rect 15788 9818 15812 9820
rect 15868 9818 15892 9820
rect 15948 9818 15954 9820
rect 15708 9766 15710 9818
rect 15890 9766 15892 9818
rect 15646 9764 15652 9766
rect 15708 9764 15732 9766
rect 15788 9764 15812 9766
rect 15868 9764 15892 9766
rect 15948 9764 15954 9766
rect 15646 9755 15954 9764
rect 15646 8732 15954 8741
rect 15646 8730 15652 8732
rect 15708 8730 15732 8732
rect 15788 8730 15812 8732
rect 15868 8730 15892 8732
rect 15948 8730 15954 8732
rect 15708 8678 15710 8730
rect 15890 8678 15892 8730
rect 15646 8676 15652 8678
rect 15708 8676 15732 8678
rect 15788 8676 15812 8678
rect 15868 8676 15892 8678
rect 15948 8676 15954 8678
rect 15646 8667 15954 8676
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15488 7546 15516 8434
rect 15646 7644 15954 7653
rect 15646 7642 15652 7644
rect 15708 7642 15732 7644
rect 15788 7642 15812 7644
rect 15868 7642 15892 7644
rect 15948 7642 15954 7644
rect 15708 7590 15710 7642
rect 15890 7590 15892 7642
rect 15646 7588 15652 7590
rect 15708 7588 15732 7590
rect 15788 7588 15812 7590
rect 15868 7588 15892 7590
rect 15948 7588 15954 7590
rect 15646 7579 15954 7588
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15488 4162 15516 5714
rect 15580 5710 15608 6598
rect 15646 6556 15954 6565
rect 15646 6554 15652 6556
rect 15708 6554 15732 6556
rect 15788 6554 15812 6556
rect 15868 6554 15892 6556
rect 15948 6554 15954 6556
rect 15708 6502 15710 6554
rect 15890 6502 15892 6554
rect 15646 6500 15652 6502
rect 15708 6500 15732 6502
rect 15788 6500 15812 6502
rect 15868 6500 15892 6502
rect 15948 6500 15954 6502
rect 15646 6491 15954 6500
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15646 5468 15954 5477
rect 15646 5466 15652 5468
rect 15708 5466 15732 5468
rect 15788 5466 15812 5468
rect 15868 5466 15892 5468
rect 15948 5466 15954 5468
rect 15708 5414 15710 5466
rect 15890 5414 15892 5466
rect 15646 5412 15652 5414
rect 15708 5412 15732 5414
rect 15788 5412 15812 5414
rect 15868 5412 15892 5414
rect 15948 5412 15954 5414
rect 15646 5403 15954 5412
rect 16040 5302 16068 8570
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 15646 4380 15954 4389
rect 15646 4378 15652 4380
rect 15708 4378 15732 4380
rect 15788 4378 15812 4380
rect 15868 4378 15892 4380
rect 15948 4378 15954 4380
rect 15708 4326 15710 4378
rect 15890 4326 15892 4378
rect 15646 4324 15652 4326
rect 15708 4324 15732 4326
rect 15788 4324 15812 4326
rect 15868 4324 15892 4326
rect 15948 4324 15954 4326
rect 15646 4315 15954 4324
rect 15488 4134 15700 4162
rect 15672 3602 15700 4134
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 15646 3292 15954 3301
rect 15646 3290 15652 3292
rect 15708 3290 15732 3292
rect 15788 3290 15812 3292
rect 15868 3290 15892 3292
rect 15948 3290 15954 3292
rect 15708 3238 15710 3290
rect 15890 3238 15892 3290
rect 15646 3236 15652 3238
rect 15708 3236 15732 3238
rect 15788 3236 15812 3238
rect 15868 3236 15892 3238
rect 15948 3236 15954 3238
rect 15646 3227 15954 3236
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 16040 2990 16068 3538
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 16132 2446 16160 9982
rect 16224 8634 16252 11630
rect 16408 10606 16436 12106
rect 16396 10600 16448 10606
rect 16396 10542 16448 10548
rect 16592 10470 16620 13194
rect 17236 12442 17264 14486
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 17144 10674 17172 11154
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 17224 10532 17276 10538
rect 17224 10474 17276 10480
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 17236 10266 17264 10474
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17328 10146 17356 16546
rect 17512 16546 17632 16574
rect 17408 16448 17460 16454
rect 17408 16390 17460 16396
rect 17420 13530 17448 16390
rect 17512 15434 17540 16546
rect 17500 15428 17552 15434
rect 17500 15370 17552 15376
rect 17696 14958 17724 17206
rect 17972 17202 18000 17478
rect 18064 17338 18092 17614
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 17960 17196 18012 17202
rect 17960 17138 18012 17144
rect 18432 16998 18460 18294
rect 18512 17604 18564 17610
rect 18512 17546 18564 17552
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18096 16892 18404 16901
rect 18096 16890 18102 16892
rect 18158 16890 18182 16892
rect 18238 16890 18262 16892
rect 18318 16890 18342 16892
rect 18398 16890 18404 16892
rect 18158 16838 18160 16890
rect 18340 16838 18342 16890
rect 18096 16836 18102 16838
rect 18158 16836 18182 16838
rect 18238 16836 18262 16838
rect 18318 16836 18342 16838
rect 18398 16836 18404 16838
rect 18096 16827 18404 16836
rect 17960 16176 18012 16182
rect 17960 16118 18012 16124
rect 17972 15162 18000 16118
rect 18524 16046 18552 17546
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18096 15804 18404 15813
rect 18096 15802 18102 15804
rect 18158 15802 18182 15804
rect 18238 15802 18262 15804
rect 18318 15802 18342 15804
rect 18398 15802 18404 15804
rect 18158 15750 18160 15802
rect 18340 15750 18342 15802
rect 18096 15748 18102 15750
rect 18158 15748 18182 15750
rect 18238 15748 18262 15750
rect 18318 15748 18342 15750
rect 18398 15748 18404 15750
rect 18096 15739 18404 15748
rect 18524 15450 18552 15982
rect 18524 15422 18644 15450
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 18524 15026 18552 15302
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18616 14958 18644 15422
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 17696 14482 17724 14894
rect 18096 14716 18404 14725
rect 18096 14714 18102 14716
rect 18158 14714 18182 14716
rect 18238 14714 18262 14716
rect 18318 14714 18342 14716
rect 18398 14714 18404 14716
rect 18158 14662 18160 14714
rect 18340 14662 18342 14714
rect 18096 14660 18102 14662
rect 18158 14660 18182 14662
rect 18238 14660 18262 14662
rect 18318 14660 18342 14662
rect 18398 14660 18404 14662
rect 18096 14651 18404 14660
rect 17684 14476 17736 14482
rect 17684 14418 17736 14424
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18432 14006 18460 14214
rect 18420 14000 18472 14006
rect 18420 13942 18472 13948
rect 18616 13870 18644 14894
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 18096 13628 18404 13637
rect 18096 13626 18102 13628
rect 18158 13626 18182 13628
rect 18238 13626 18262 13628
rect 18318 13626 18342 13628
rect 18398 13626 18404 13628
rect 18158 13574 18160 13626
rect 18340 13574 18342 13626
rect 18096 13572 18102 13574
rect 18158 13572 18182 13574
rect 18238 13572 18262 13574
rect 18318 13572 18342 13574
rect 18398 13572 18404 13574
rect 18096 13563 18404 13572
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17420 13326 17448 13466
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 18064 12850 18092 13126
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18096 12540 18404 12549
rect 18096 12538 18102 12540
rect 18158 12538 18182 12540
rect 18238 12538 18262 12540
rect 18318 12538 18342 12540
rect 18398 12538 18404 12540
rect 18158 12486 18160 12538
rect 18340 12486 18342 12538
rect 18096 12484 18102 12486
rect 18158 12484 18182 12486
rect 18238 12484 18262 12486
rect 18318 12484 18342 12486
rect 18398 12484 18404 12486
rect 18096 12475 18404 12484
rect 17592 12368 17644 12374
rect 17592 12310 17644 12316
rect 17604 10810 17632 12310
rect 18432 12238 18460 12582
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 18096 11452 18404 11461
rect 18096 11450 18102 11452
rect 18158 11450 18182 11452
rect 18238 11450 18262 11452
rect 18318 11450 18342 11452
rect 18398 11450 18404 11452
rect 18158 11398 18160 11450
rect 18340 11398 18342 11450
rect 18096 11396 18102 11398
rect 18158 11396 18182 11398
rect 18238 11396 18262 11398
rect 18318 11396 18342 11398
rect 18398 11396 18404 11398
rect 18096 11387 18404 11396
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 18616 10606 18644 13806
rect 18984 13258 19012 20810
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19248 15360 19300 15366
rect 19248 15302 19300 15308
rect 19352 15314 19380 15642
rect 19444 15434 19472 20742
rect 19616 20528 19668 20534
rect 19616 20470 19668 20476
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19432 15428 19484 15434
rect 19432 15370 19484 15376
rect 19260 15065 19288 15302
rect 19352 15286 19472 15314
rect 19246 15056 19302 15065
rect 19246 14991 19302 15000
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18892 11830 18920 12038
rect 19444 11830 19472 15286
rect 18880 11824 18932 11830
rect 18880 11766 18932 11772
rect 19432 11824 19484 11830
rect 19432 11766 19484 11772
rect 19444 10742 19472 11766
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 17408 10600 17460 10606
rect 17408 10542 17460 10548
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 17144 10118 17356 10146
rect 17420 10130 17448 10542
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17408 10124 17460 10130
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16304 8356 16356 8362
rect 16304 8298 16356 8304
rect 16316 7954 16344 8298
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16592 7410 16620 7890
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16224 5778 16252 6054
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 16224 5642 16252 5714
rect 16212 5636 16264 5642
rect 16212 5578 16264 5584
rect 16224 3466 16252 5578
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 16224 3194 16252 3402
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 17144 3058 17172 10118
rect 17408 10066 17460 10072
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17236 7546 17264 8434
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 17328 7410 17356 8230
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 17512 6914 17540 10406
rect 18096 10364 18404 10373
rect 18096 10362 18102 10364
rect 18158 10362 18182 10364
rect 18238 10362 18262 10364
rect 18318 10362 18342 10364
rect 18398 10362 18404 10364
rect 18158 10310 18160 10362
rect 18340 10310 18342 10362
rect 18096 10308 18102 10310
rect 18158 10308 18182 10310
rect 18238 10308 18262 10310
rect 18318 10308 18342 10310
rect 18398 10308 18404 10310
rect 18096 10299 18404 10308
rect 17592 10192 17644 10198
rect 17592 10134 17644 10140
rect 17420 6886 17540 6914
rect 17604 6914 17632 10134
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18096 9276 18404 9285
rect 18096 9274 18102 9276
rect 18158 9274 18182 9276
rect 18238 9274 18262 9276
rect 18318 9274 18342 9276
rect 18398 9274 18404 9276
rect 18158 9222 18160 9274
rect 18340 9222 18342 9274
rect 18096 9220 18102 9222
rect 18158 9220 18182 9222
rect 18238 9220 18262 9222
rect 18318 9220 18342 9222
rect 18398 9220 18404 9222
rect 18096 9211 18404 9220
rect 18524 8566 18552 9862
rect 18420 8560 18472 8566
rect 18420 8502 18472 8508
rect 18512 8560 18564 8566
rect 18512 8502 18564 8508
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17696 7546 17724 8366
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17604 6886 17724 6914
rect 17420 6458 17448 6886
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17420 6118 17448 6394
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17696 5642 17724 6886
rect 17880 6866 17908 8434
rect 18432 8378 18460 8502
rect 18616 8430 18644 10542
rect 19444 8566 19472 10678
rect 19432 8560 19484 8566
rect 19432 8502 19484 8508
rect 18604 8424 18656 8430
rect 17960 8356 18012 8362
rect 18432 8350 18552 8378
rect 18604 8366 18656 8372
rect 17960 8298 18012 8304
rect 17972 7410 18000 8298
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18096 8188 18404 8197
rect 18096 8186 18102 8188
rect 18158 8186 18182 8188
rect 18238 8186 18262 8188
rect 18318 8186 18342 8188
rect 18398 8186 18404 8188
rect 18158 8134 18160 8186
rect 18340 8134 18342 8186
rect 18096 8132 18102 8134
rect 18158 8132 18182 8134
rect 18238 8132 18262 8134
rect 18318 8132 18342 8134
rect 18398 8132 18404 8134
rect 18096 8123 18404 8132
rect 18432 7886 18460 8230
rect 18524 8090 18552 8350
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18616 7970 18644 8366
rect 18524 7942 18644 7970
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 18420 7336 18472 7342
rect 18420 7278 18472 7284
rect 18096 7100 18404 7109
rect 18096 7098 18102 7100
rect 18158 7098 18182 7100
rect 18238 7098 18262 7100
rect 18318 7098 18342 7100
rect 18398 7098 18404 7100
rect 18158 7046 18160 7098
rect 18340 7046 18342 7098
rect 18096 7044 18102 7046
rect 18158 7044 18182 7046
rect 18238 7044 18262 7046
rect 18318 7044 18342 7046
rect 18398 7044 18404 7046
rect 18096 7035 18404 7044
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 18432 6322 18460 7278
rect 18524 6322 18552 7942
rect 18604 7812 18656 7818
rect 18604 7754 18656 7760
rect 18616 7410 18644 7754
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 19444 6866 19472 8502
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19444 6390 19472 6802
rect 19432 6384 19484 6390
rect 19432 6326 19484 6332
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17788 5710 17816 6054
rect 18096 6012 18404 6021
rect 18096 6010 18102 6012
rect 18158 6010 18182 6012
rect 18238 6010 18262 6012
rect 18318 6010 18342 6012
rect 18398 6010 18404 6012
rect 18158 5958 18160 6010
rect 18340 5958 18342 6010
rect 18096 5956 18102 5958
rect 18158 5956 18182 5958
rect 18238 5956 18262 5958
rect 18318 5956 18342 5958
rect 18398 5956 18404 5958
rect 18096 5947 18404 5956
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 17684 5636 17736 5642
rect 17684 5578 17736 5584
rect 17592 5568 17644 5574
rect 17592 5510 17644 5516
rect 17604 4010 17632 5510
rect 18432 5370 18460 5646
rect 18420 5364 18472 5370
rect 18420 5306 18472 5312
rect 18524 5234 18552 6258
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 18892 5914 18920 6190
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 19444 5386 19472 6326
rect 19352 5358 19472 5386
rect 19352 5302 19380 5358
rect 19248 5296 19300 5302
rect 19340 5296 19392 5302
rect 19300 5244 19340 5250
rect 19248 5238 19392 5244
rect 18512 5228 18564 5234
rect 19260 5222 19380 5238
rect 18512 5170 18564 5176
rect 18096 4924 18404 4933
rect 18096 4922 18102 4924
rect 18158 4922 18182 4924
rect 18238 4922 18262 4924
rect 18318 4922 18342 4924
rect 18398 4922 18404 4924
rect 18158 4870 18160 4922
rect 18340 4870 18342 4922
rect 18096 4868 18102 4870
rect 18158 4868 18182 4870
rect 18238 4868 18262 4870
rect 18318 4868 18342 4870
rect 18398 4868 18404 4870
rect 18096 4859 18404 4868
rect 18524 4146 18552 5170
rect 18788 5160 18840 5166
rect 18788 5102 18840 5108
rect 18800 4826 18828 5102
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 19352 4214 19380 5222
rect 19340 4208 19392 4214
rect 19340 4150 19392 4156
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 17592 4004 17644 4010
rect 17592 3946 17644 3952
rect 18096 3836 18404 3845
rect 18096 3834 18102 3836
rect 18158 3834 18182 3836
rect 18238 3834 18262 3836
rect 18318 3834 18342 3836
rect 18398 3834 18404 3836
rect 18158 3782 18160 3834
rect 18340 3782 18342 3834
rect 18096 3780 18102 3782
rect 18158 3780 18182 3782
rect 18238 3780 18262 3782
rect 18318 3780 18342 3782
rect 18398 3780 18404 3782
rect 18096 3771 18404 3780
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17420 2446 17448 3334
rect 18972 2848 19024 2854
rect 18972 2790 19024 2796
rect 18096 2748 18404 2757
rect 18096 2746 18102 2748
rect 18158 2746 18182 2748
rect 18238 2746 18262 2748
rect 18318 2746 18342 2748
rect 18398 2746 18404 2748
rect 18158 2694 18160 2746
rect 18340 2694 18342 2746
rect 18096 2692 18102 2694
rect 18158 2692 18182 2694
rect 18238 2692 18262 2694
rect 18318 2692 18342 2694
rect 18398 2692 18404 2694
rect 18096 2683 18404 2692
rect 18984 2446 19012 2790
rect 19536 2446 19564 18022
rect 19628 17882 19656 20470
rect 19720 19514 19748 21490
rect 21192 21146 21220 23224
rect 21180 21140 21232 21146
rect 21180 21082 21232 21088
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 20260 20868 20312 20874
rect 20260 20810 20312 20816
rect 19708 19508 19760 19514
rect 19708 19450 19760 19456
rect 20076 18760 20128 18766
rect 20076 18702 20128 18708
rect 20088 17882 20116 18702
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 19628 17270 19656 17818
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 19616 17264 19668 17270
rect 19616 17206 19668 17212
rect 19892 16720 19944 16726
rect 19892 16662 19944 16668
rect 19904 16114 19932 16662
rect 19984 16516 20036 16522
rect 19984 16458 20036 16464
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 19800 15496 19852 15502
rect 19800 15438 19852 15444
rect 19812 15162 19840 15438
rect 19800 15156 19852 15162
rect 19800 15098 19852 15104
rect 19904 15094 19932 16050
rect 19996 15706 20024 16458
rect 20088 16250 20116 17614
rect 20180 16522 20208 20810
rect 20272 20602 20300 20810
rect 20545 20700 20853 20709
rect 20545 20698 20551 20700
rect 20607 20698 20631 20700
rect 20687 20698 20711 20700
rect 20767 20698 20791 20700
rect 20847 20698 20853 20700
rect 20607 20646 20609 20698
rect 20789 20646 20791 20698
rect 20545 20644 20551 20646
rect 20607 20644 20631 20646
rect 20687 20644 20711 20646
rect 20767 20644 20791 20646
rect 20847 20644 20853 20646
rect 20545 20635 20853 20644
rect 20260 20596 20312 20602
rect 20260 20538 20312 20544
rect 20350 19952 20406 19961
rect 20350 19887 20406 19896
rect 20364 19854 20392 19887
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20545 19612 20853 19621
rect 20545 19610 20551 19612
rect 20607 19610 20631 19612
rect 20687 19610 20711 19612
rect 20767 19610 20791 19612
rect 20847 19610 20853 19612
rect 20607 19558 20609 19610
rect 20789 19558 20791 19610
rect 20545 19556 20551 19558
rect 20607 19556 20631 19558
rect 20687 19556 20711 19558
rect 20767 19556 20791 19558
rect 20847 19556 20853 19558
rect 20545 19547 20853 19556
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20272 18329 20300 18566
rect 20545 18524 20853 18533
rect 20545 18522 20551 18524
rect 20607 18522 20631 18524
rect 20687 18522 20711 18524
rect 20767 18522 20791 18524
rect 20847 18522 20853 18524
rect 20607 18470 20609 18522
rect 20789 18470 20791 18522
rect 20545 18468 20551 18470
rect 20607 18468 20631 18470
rect 20687 18468 20711 18470
rect 20767 18468 20791 18470
rect 20847 18468 20853 18470
rect 20545 18459 20853 18468
rect 20258 18320 20314 18329
rect 20258 18255 20314 18264
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 20272 16697 20300 17478
rect 20545 17436 20853 17445
rect 20545 17434 20551 17436
rect 20607 17434 20631 17436
rect 20687 17434 20711 17436
rect 20767 17434 20791 17436
rect 20847 17434 20853 17436
rect 20607 17382 20609 17434
rect 20789 17382 20791 17434
rect 20545 17380 20551 17382
rect 20607 17380 20631 17382
rect 20687 17380 20711 17382
rect 20767 17380 20791 17382
rect 20847 17380 20853 17382
rect 20545 17371 20853 17380
rect 20444 16992 20496 16998
rect 20444 16934 20496 16940
rect 20258 16688 20314 16697
rect 20258 16623 20314 16632
rect 20168 16516 20220 16522
rect 20168 16458 20220 16464
rect 20076 16244 20128 16250
rect 20076 16186 20128 16192
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 19892 15088 19944 15094
rect 19892 15030 19944 15036
rect 19904 14006 19932 15030
rect 19892 14000 19944 14006
rect 19892 13942 19944 13948
rect 20352 13728 20404 13734
rect 20352 13670 20404 13676
rect 20168 13456 20220 13462
rect 20166 13424 20168 13433
rect 20220 13424 20222 13433
rect 20166 13359 20222 13368
rect 20364 13326 20392 13670
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 20352 12232 20404 12238
rect 20352 12174 20404 12180
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 20180 11801 20208 12038
rect 20364 11898 20392 12174
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20166 11792 20222 11801
rect 20166 11727 20222 11736
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20168 10192 20220 10198
rect 20166 10160 20168 10169
rect 20220 10160 20222 10169
rect 20166 10095 20222 10104
rect 20364 10062 20392 10406
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 20180 8537 20208 8774
rect 20364 8634 20392 8910
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20166 8528 20222 8537
rect 20166 8463 20222 8472
rect 20166 6896 20222 6905
rect 20166 6831 20222 6840
rect 20180 6662 20208 6831
rect 20352 6792 20404 6798
rect 20352 6734 20404 6740
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20364 6458 20392 6734
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20272 5273 20300 5510
rect 20258 5264 20314 5273
rect 20258 5199 20314 5208
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 20088 3534 20116 4966
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 20260 3664 20312 3670
rect 20258 3632 20260 3641
rect 20312 3632 20314 3641
rect 20258 3567 20314 3576
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 20364 3058 20392 3878
rect 20352 3052 20404 3058
rect 20352 2994 20404 3000
rect 20168 2848 20220 2854
rect 20168 2790 20220 2796
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 18972 2440 19024 2446
rect 18972 2382 19024 2388
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 13452 2304 13504 2310
rect 13452 2246 13504 2252
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 19892 2304 19944 2310
rect 19892 2246 19944 2252
rect 10747 2204 11055 2213
rect 10747 2202 10753 2204
rect 10809 2202 10833 2204
rect 10889 2202 10913 2204
rect 10969 2202 10993 2204
rect 11049 2202 11055 2204
rect 10809 2150 10811 2202
rect 10991 2150 10993 2202
rect 10747 2148 10753 2150
rect 10809 2148 10833 2150
rect 10889 2148 10913 2150
rect 10969 2148 10993 2150
rect 11049 2148 11055 2150
rect 10747 2139 11055 2148
rect 10796 870 10916 898
rect 10796 762 10824 870
rect 10888 800 10916 870
rect 12176 800 12204 2246
rect 13464 800 13492 2246
rect 14752 800 14780 2246
rect 15646 2204 15954 2213
rect 15646 2202 15652 2204
rect 15708 2202 15732 2204
rect 15788 2202 15812 2204
rect 15868 2202 15892 2204
rect 15948 2202 15954 2204
rect 15708 2150 15710 2202
rect 15890 2150 15892 2202
rect 15646 2148 15652 2150
rect 15708 2148 15732 2150
rect 15788 2148 15812 2150
rect 15868 2148 15892 2150
rect 15948 2148 15954 2150
rect 15646 2139 15954 2148
rect 16040 800 16068 2246
rect 17328 800 17356 2246
rect 18616 800 18644 2246
rect 19904 800 19932 2246
rect 20180 2009 20208 2790
rect 20456 2446 20484 16934
rect 20545 16348 20853 16357
rect 20545 16346 20551 16348
rect 20607 16346 20631 16348
rect 20687 16346 20711 16348
rect 20767 16346 20791 16348
rect 20847 16346 20853 16348
rect 20607 16294 20609 16346
rect 20789 16294 20791 16346
rect 20545 16292 20551 16294
rect 20607 16292 20631 16294
rect 20687 16292 20711 16294
rect 20767 16292 20791 16294
rect 20847 16292 20853 16294
rect 20545 16283 20853 16292
rect 20545 15260 20853 15269
rect 20545 15258 20551 15260
rect 20607 15258 20631 15260
rect 20687 15258 20711 15260
rect 20767 15258 20791 15260
rect 20847 15258 20853 15260
rect 20607 15206 20609 15258
rect 20789 15206 20791 15258
rect 20545 15204 20551 15206
rect 20607 15204 20631 15206
rect 20687 15204 20711 15206
rect 20767 15204 20791 15206
rect 20847 15204 20853 15206
rect 20545 15195 20853 15204
rect 20545 14172 20853 14181
rect 20545 14170 20551 14172
rect 20607 14170 20631 14172
rect 20687 14170 20711 14172
rect 20767 14170 20791 14172
rect 20847 14170 20853 14172
rect 20607 14118 20609 14170
rect 20789 14118 20791 14170
rect 20545 14116 20551 14118
rect 20607 14116 20631 14118
rect 20687 14116 20711 14118
rect 20767 14116 20791 14118
rect 20847 14116 20853 14118
rect 20545 14107 20853 14116
rect 20545 13084 20853 13093
rect 20545 13082 20551 13084
rect 20607 13082 20631 13084
rect 20687 13082 20711 13084
rect 20767 13082 20791 13084
rect 20847 13082 20853 13084
rect 20607 13030 20609 13082
rect 20789 13030 20791 13082
rect 20545 13028 20551 13030
rect 20607 13028 20631 13030
rect 20687 13028 20711 13030
rect 20767 13028 20791 13030
rect 20847 13028 20853 13030
rect 20545 13019 20853 13028
rect 20545 11996 20853 12005
rect 20545 11994 20551 11996
rect 20607 11994 20631 11996
rect 20687 11994 20711 11996
rect 20767 11994 20791 11996
rect 20847 11994 20853 11996
rect 20607 11942 20609 11994
rect 20789 11942 20791 11994
rect 20545 11940 20551 11942
rect 20607 11940 20631 11942
rect 20687 11940 20711 11942
rect 20767 11940 20791 11942
rect 20847 11940 20853 11942
rect 20545 11931 20853 11940
rect 20545 10908 20853 10917
rect 20545 10906 20551 10908
rect 20607 10906 20631 10908
rect 20687 10906 20711 10908
rect 20767 10906 20791 10908
rect 20847 10906 20853 10908
rect 20607 10854 20609 10906
rect 20789 10854 20791 10906
rect 20545 10852 20551 10854
rect 20607 10852 20631 10854
rect 20687 10852 20711 10854
rect 20767 10852 20791 10854
rect 20847 10852 20853 10854
rect 20545 10843 20853 10852
rect 20545 9820 20853 9829
rect 20545 9818 20551 9820
rect 20607 9818 20631 9820
rect 20687 9818 20711 9820
rect 20767 9818 20791 9820
rect 20847 9818 20853 9820
rect 20607 9766 20609 9818
rect 20789 9766 20791 9818
rect 20545 9764 20551 9766
rect 20607 9764 20631 9766
rect 20687 9764 20711 9766
rect 20767 9764 20791 9766
rect 20847 9764 20853 9766
rect 20545 9755 20853 9764
rect 20545 8732 20853 8741
rect 20545 8730 20551 8732
rect 20607 8730 20631 8732
rect 20687 8730 20711 8732
rect 20767 8730 20791 8732
rect 20847 8730 20853 8732
rect 20607 8678 20609 8730
rect 20789 8678 20791 8730
rect 20545 8676 20551 8678
rect 20607 8676 20631 8678
rect 20687 8676 20711 8678
rect 20767 8676 20791 8678
rect 20847 8676 20853 8678
rect 20545 8667 20853 8676
rect 20545 7644 20853 7653
rect 20545 7642 20551 7644
rect 20607 7642 20631 7644
rect 20687 7642 20711 7644
rect 20767 7642 20791 7644
rect 20847 7642 20853 7644
rect 20607 7590 20609 7642
rect 20789 7590 20791 7642
rect 20545 7588 20551 7590
rect 20607 7588 20631 7590
rect 20687 7588 20711 7590
rect 20767 7588 20791 7590
rect 20847 7588 20853 7590
rect 20545 7579 20853 7588
rect 20545 6556 20853 6565
rect 20545 6554 20551 6556
rect 20607 6554 20631 6556
rect 20687 6554 20711 6556
rect 20767 6554 20791 6556
rect 20847 6554 20853 6556
rect 20607 6502 20609 6554
rect 20789 6502 20791 6554
rect 20545 6500 20551 6502
rect 20607 6500 20631 6502
rect 20687 6500 20711 6502
rect 20767 6500 20791 6502
rect 20847 6500 20853 6502
rect 20545 6491 20853 6500
rect 20545 5468 20853 5477
rect 20545 5466 20551 5468
rect 20607 5466 20631 5468
rect 20687 5466 20711 5468
rect 20767 5466 20791 5468
rect 20847 5466 20853 5468
rect 20607 5414 20609 5466
rect 20789 5414 20791 5466
rect 20545 5412 20551 5414
rect 20607 5412 20631 5414
rect 20687 5412 20711 5414
rect 20767 5412 20791 5414
rect 20847 5412 20853 5414
rect 20545 5403 20853 5412
rect 20545 4380 20853 4389
rect 20545 4378 20551 4380
rect 20607 4378 20631 4380
rect 20687 4378 20711 4380
rect 20767 4378 20791 4380
rect 20847 4378 20853 4380
rect 20607 4326 20609 4378
rect 20789 4326 20791 4378
rect 20545 4324 20551 4326
rect 20607 4324 20631 4326
rect 20687 4324 20711 4326
rect 20767 4324 20791 4326
rect 20847 4324 20853 4326
rect 20545 4315 20853 4324
rect 20545 3292 20853 3301
rect 20545 3290 20551 3292
rect 20607 3290 20631 3292
rect 20687 3290 20711 3292
rect 20767 3290 20791 3292
rect 20847 3290 20853 3292
rect 20607 3238 20609 3290
rect 20789 3238 20791 3290
rect 20545 3236 20551 3238
rect 20607 3236 20631 3238
rect 20687 3236 20711 3238
rect 20767 3236 20791 3238
rect 20847 3236 20853 3238
rect 20545 3227 20853 3236
rect 20444 2440 20496 2446
rect 20444 2382 20496 2388
rect 21180 2304 21232 2310
rect 21180 2246 21232 2252
rect 20545 2204 20853 2213
rect 20545 2202 20551 2204
rect 20607 2202 20631 2204
rect 20687 2202 20711 2204
rect 20767 2202 20791 2204
rect 20847 2202 20853 2204
rect 20607 2150 20609 2202
rect 20789 2150 20791 2202
rect 20545 2148 20551 2150
rect 20607 2148 20631 2150
rect 20687 2148 20711 2150
rect 20767 2148 20791 2150
rect 20847 2148 20853 2150
rect 20545 2139 20853 2148
rect 20166 2000 20222 2009
rect 20166 1935 20222 1944
rect 21192 800 21220 2246
rect 10612 734 10824 762
rect 10874 0 10930 800
rect 12162 0 12218 800
rect 13450 0 13506 800
rect 14738 0 14794 800
rect 16026 0 16082 800
rect 17314 0 17370 800
rect 18602 0 18658 800
rect 19890 0 19946 800
rect 21178 0 21234 800
<< via2 >>
rect 5854 21786 5910 21788
rect 5934 21786 5990 21788
rect 6014 21786 6070 21788
rect 6094 21786 6150 21788
rect 5854 21734 5900 21786
rect 5900 21734 5910 21786
rect 5934 21734 5964 21786
rect 5964 21734 5976 21786
rect 5976 21734 5990 21786
rect 6014 21734 6028 21786
rect 6028 21734 6040 21786
rect 6040 21734 6070 21786
rect 6094 21734 6104 21786
rect 6104 21734 6150 21786
rect 5854 21732 5910 21734
rect 5934 21732 5990 21734
rect 6014 21732 6070 21734
rect 6094 21732 6150 21734
rect 10753 21786 10809 21788
rect 10833 21786 10889 21788
rect 10913 21786 10969 21788
rect 10993 21786 11049 21788
rect 10753 21734 10799 21786
rect 10799 21734 10809 21786
rect 10833 21734 10863 21786
rect 10863 21734 10875 21786
rect 10875 21734 10889 21786
rect 10913 21734 10927 21786
rect 10927 21734 10939 21786
rect 10939 21734 10969 21786
rect 10993 21734 11003 21786
rect 11003 21734 11049 21786
rect 10753 21732 10809 21734
rect 10833 21732 10889 21734
rect 10913 21732 10969 21734
rect 10993 21732 11049 21734
rect 15652 21786 15708 21788
rect 15732 21786 15788 21788
rect 15812 21786 15868 21788
rect 15892 21786 15948 21788
rect 15652 21734 15698 21786
rect 15698 21734 15708 21786
rect 15732 21734 15762 21786
rect 15762 21734 15774 21786
rect 15774 21734 15788 21786
rect 15812 21734 15826 21786
rect 15826 21734 15838 21786
rect 15838 21734 15868 21786
rect 15892 21734 15902 21786
rect 15902 21734 15948 21786
rect 15652 21732 15708 21734
rect 15732 21732 15788 21734
rect 15812 21732 15868 21734
rect 15892 21732 15948 21734
rect 20551 21786 20607 21788
rect 20631 21786 20687 21788
rect 20711 21786 20767 21788
rect 20791 21786 20847 21788
rect 20551 21734 20597 21786
rect 20597 21734 20607 21786
rect 20631 21734 20661 21786
rect 20661 21734 20673 21786
rect 20673 21734 20687 21786
rect 20711 21734 20725 21786
rect 20725 21734 20737 21786
rect 20737 21734 20767 21786
rect 20791 21734 20801 21786
rect 20801 21734 20847 21786
rect 20551 21732 20607 21734
rect 20631 21732 20687 21734
rect 20711 21732 20767 21734
rect 20791 21732 20847 21734
rect 19614 21528 19670 21584
rect 1306 21256 1362 21312
rect 1398 13640 1454 13696
rect 846 10004 848 10024
rect 848 10004 900 10024
rect 900 10004 902 10024
rect 846 9968 902 10004
rect 3405 21242 3461 21244
rect 3485 21242 3541 21244
rect 3565 21242 3621 21244
rect 3645 21242 3701 21244
rect 3405 21190 3451 21242
rect 3451 21190 3461 21242
rect 3485 21190 3515 21242
rect 3515 21190 3527 21242
rect 3527 21190 3541 21242
rect 3565 21190 3579 21242
rect 3579 21190 3591 21242
rect 3591 21190 3621 21242
rect 3645 21190 3655 21242
rect 3655 21190 3701 21242
rect 3405 21188 3461 21190
rect 3485 21188 3541 21190
rect 3565 21188 3621 21190
rect 3645 21188 3701 21190
rect 3405 20154 3461 20156
rect 3485 20154 3541 20156
rect 3565 20154 3621 20156
rect 3645 20154 3701 20156
rect 3405 20102 3451 20154
rect 3451 20102 3461 20154
rect 3485 20102 3515 20154
rect 3515 20102 3527 20154
rect 3527 20102 3541 20154
rect 3565 20102 3579 20154
rect 3579 20102 3591 20154
rect 3591 20102 3621 20154
rect 3645 20102 3655 20154
rect 3655 20102 3701 20154
rect 3405 20100 3461 20102
rect 3485 20100 3541 20102
rect 3565 20100 3621 20102
rect 3645 20100 3701 20102
rect 3405 19066 3461 19068
rect 3485 19066 3541 19068
rect 3565 19066 3621 19068
rect 3645 19066 3701 19068
rect 3405 19014 3451 19066
rect 3451 19014 3461 19066
rect 3485 19014 3515 19066
rect 3515 19014 3527 19066
rect 3527 19014 3541 19066
rect 3565 19014 3579 19066
rect 3579 19014 3591 19066
rect 3591 19014 3621 19066
rect 3645 19014 3655 19066
rect 3655 19014 3701 19066
rect 3405 19012 3461 19014
rect 3485 19012 3541 19014
rect 3565 19012 3621 19014
rect 3645 19012 3701 19014
rect 3405 17978 3461 17980
rect 3485 17978 3541 17980
rect 3565 17978 3621 17980
rect 3645 17978 3701 17980
rect 3405 17926 3451 17978
rect 3451 17926 3461 17978
rect 3485 17926 3515 17978
rect 3515 17926 3527 17978
rect 3527 17926 3541 17978
rect 3565 17926 3579 17978
rect 3579 17926 3591 17978
rect 3591 17926 3621 17978
rect 3645 17926 3655 17978
rect 3655 17926 3701 17978
rect 3405 17924 3461 17926
rect 3485 17924 3541 17926
rect 3565 17924 3621 17926
rect 3645 17924 3701 17926
rect 3405 16890 3461 16892
rect 3485 16890 3541 16892
rect 3565 16890 3621 16892
rect 3645 16890 3701 16892
rect 3405 16838 3451 16890
rect 3451 16838 3461 16890
rect 3485 16838 3515 16890
rect 3515 16838 3527 16890
rect 3527 16838 3541 16890
rect 3565 16838 3579 16890
rect 3579 16838 3591 16890
rect 3591 16838 3621 16890
rect 3645 16838 3655 16890
rect 3655 16838 3701 16890
rect 3405 16836 3461 16838
rect 3485 16836 3541 16838
rect 3565 16836 3621 16838
rect 3645 16836 3701 16838
rect 3405 15802 3461 15804
rect 3485 15802 3541 15804
rect 3565 15802 3621 15804
rect 3645 15802 3701 15804
rect 3405 15750 3451 15802
rect 3451 15750 3461 15802
rect 3485 15750 3515 15802
rect 3515 15750 3527 15802
rect 3527 15750 3541 15802
rect 3565 15750 3579 15802
rect 3579 15750 3591 15802
rect 3591 15750 3621 15802
rect 3645 15750 3655 15802
rect 3655 15750 3701 15802
rect 3405 15748 3461 15750
rect 3485 15748 3541 15750
rect 3565 15748 3621 15750
rect 3645 15748 3701 15750
rect 3405 14714 3461 14716
rect 3485 14714 3541 14716
rect 3565 14714 3621 14716
rect 3645 14714 3701 14716
rect 3405 14662 3451 14714
rect 3451 14662 3461 14714
rect 3485 14662 3515 14714
rect 3515 14662 3527 14714
rect 3527 14662 3541 14714
rect 3565 14662 3579 14714
rect 3579 14662 3591 14714
rect 3591 14662 3621 14714
rect 3645 14662 3655 14714
rect 3655 14662 3701 14714
rect 3405 14660 3461 14662
rect 3485 14660 3541 14662
rect 3565 14660 3621 14662
rect 3645 14660 3701 14662
rect 3405 13626 3461 13628
rect 3485 13626 3541 13628
rect 3565 13626 3621 13628
rect 3645 13626 3701 13628
rect 3405 13574 3451 13626
rect 3451 13574 3461 13626
rect 3485 13574 3515 13626
rect 3515 13574 3527 13626
rect 3527 13574 3541 13626
rect 3565 13574 3579 13626
rect 3579 13574 3591 13626
rect 3591 13574 3621 13626
rect 3645 13574 3655 13626
rect 3655 13574 3701 13626
rect 3405 13572 3461 13574
rect 3485 13572 3541 13574
rect 3565 13572 3621 13574
rect 3645 13572 3701 13574
rect 3405 12538 3461 12540
rect 3485 12538 3541 12540
rect 3565 12538 3621 12540
rect 3645 12538 3701 12540
rect 3405 12486 3451 12538
rect 3451 12486 3461 12538
rect 3485 12486 3515 12538
rect 3515 12486 3527 12538
rect 3527 12486 3541 12538
rect 3565 12486 3579 12538
rect 3579 12486 3591 12538
rect 3591 12486 3621 12538
rect 3645 12486 3655 12538
rect 3655 12486 3701 12538
rect 3405 12484 3461 12486
rect 3485 12484 3541 12486
rect 3565 12484 3621 12486
rect 3645 12484 3701 12486
rect 3405 11450 3461 11452
rect 3485 11450 3541 11452
rect 3565 11450 3621 11452
rect 3645 11450 3701 11452
rect 3405 11398 3451 11450
rect 3451 11398 3461 11450
rect 3485 11398 3515 11450
rect 3515 11398 3527 11450
rect 3527 11398 3541 11450
rect 3565 11398 3579 11450
rect 3579 11398 3591 11450
rect 3591 11398 3621 11450
rect 3645 11398 3655 11450
rect 3655 11398 3701 11450
rect 3405 11396 3461 11398
rect 3485 11396 3541 11398
rect 3565 11396 3621 11398
rect 3645 11396 3701 11398
rect 3405 10362 3461 10364
rect 3485 10362 3541 10364
rect 3565 10362 3621 10364
rect 3645 10362 3701 10364
rect 3405 10310 3451 10362
rect 3451 10310 3461 10362
rect 3485 10310 3515 10362
rect 3515 10310 3527 10362
rect 3527 10310 3541 10362
rect 3565 10310 3579 10362
rect 3579 10310 3591 10362
rect 3591 10310 3621 10362
rect 3645 10310 3655 10362
rect 3655 10310 3701 10362
rect 3405 10308 3461 10310
rect 3485 10308 3541 10310
rect 3565 10308 3621 10310
rect 3645 10308 3701 10310
rect 3405 9274 3461 9276
rect 3485 9274 3541 9276
rect 3565 9274 3621 9276
rect 3645 9274 3701 9276
rect 3405 9222 3451 9274
rect 3451 9222 3461 9274
rect 3485 9222 3515 9274
rect 3515 9222 3527 9274
rect 3527 9222 3541 9274
rect 3565 9222 3579 9274
rect 3579 9222 3591 9274
rect 3591 9222 3621 9274
rect 3645 9222 3655 9274
rect 3655 9222 3701 9274
rect 3405 9220 3461 9222
rect 3485 9220 3541 9222
rect 3565 9220 3621 9222
rect 3645 9220 3701 9222
rect 3405 8186 3461 8188
rect 3485 8186 3541 8188
rect 3565 8186 3621 8188
rect 3645 8186 3701 8188
rect 3405 8134 3451 8186
rect 3451 8134 3461 8186
rect 3485 8134 3515 8186
rect 3515 8134 3527 8186
rect 3527 8134 3541 8186
rect 3565 8134 3579 8186
rect 3579 8134 3591 8186
rect 3591 8134 3621 8186
rect 3645 8134 3655 8186
rect 3655 8134 3701 8186
rect 3405 8132 3461 8134
rect 3485 8132 3541 8134
rect 3565 8132 3621 8134
rect 3645 8132 3701 8134
rect 3405 7098 3461 7100
rect 3485 7098 3541 7100
rect 3565 7098 3621 7100
rect 3645 7098 3701 7100
rect 3405 7046 3451 7098
rect 3451 7046 3461 7098
rect 3485 7046 3515 7098
rect 3515 7046 3527 7098
rect 3527 7046 3541 7098
rect 3565 7046 3579 7098
rect 3579 7046 3591 7098
rect 3591 7046 3621 7098
rect 3645 7046 3655 7098
rect 3655 7046 3701 7098
rect 3405 7044 3461 7046
rect 3485 7044 3541 7046
rect 3565 7044 3621 7046
rect 3645 7044 3701 7046
rect 3405 6010 3461 6012
rect 3485 6010 3541 6012
rect 3565 6010 3621 6012
rect 3645 6010 3701 6012
rect 3405 5958 3451 6010
rect 3451 5958 3461 6010
rect 3485 5958 3515 6010
rect 3515 5958 3527 6010
rect 3527 5958 3541 6010
rect 3565 5958 3579 6010
rect 3579 5958 3591 6010
rect 3591 5958 3621 6010
rect 3645 5958 3655 6010
rect 3655 5958 3701 6010
rect 3405 5956 3461 5958
rect 3485 5956 3541 5958
rect 3565 5956 3621 5958
rect 3645 5956 3701 5958
rect 3405 4922 3461 4924
rect 3485 4922 3541 4924
rect 3565 4922 3621 4924
rect 3645 4922 3701 4924
rect 3405 4870 3451 4922
rect 3451 4870 3461 4922
rect 3485 4870 3515 4922
rect 3515 4870 3527 4922
rect 3527 4870 3541 4922
rect 3565 4870 3579 4922
rect 3579 4870 3591 4922
rect 3591 4870 3621 4922
rect 3645 4870 3655 4922
rect 3655 4870 3701 4922
rect 3405 4868 3461 4870
rect 3485 4868 3541 4870
rect 3565 4868 3621 4870
rect 3645 4868 3701 4870
rect 3405 3834 3461 3836
rect 3485 3834 3541 3836
rect 3565 3834 3621 3836
rect 3645 3834 3701 3836
rect 3405 3782 3451 3834
rect 3451 3782 3461 3834
rect 3485 3782 3515 3834
rect 3515 3782 3527 3834
rect 3527 3782 3541 3834
rect 3565 3782 3579 3834
rect 3579 3782 3591 3834
rect 3591 3782 3621 3834
rect 3645 3782 3655 3834
rect 3655 3782 3701 3834
rect 3405 3780 3461 3782
rect 3485 3780 3541 3782
rect 3565 3780 3621 3782
rect 3645 3780 3701 3782
rect 3405 2746 3461 2748
rect 3485 2746 3541 2748
rect 3565 2746 3621 2748
rect 3645 2746 3701 2748
rect 3405 2694 3451 2746
rect 3451 2694 3461 2746
rect 3485 2694 3515 2746
rect 3515 2694 3527 2746
rect 3527 2694 3541 2746
rect 3565 2694 3579 2746
rect 3579 2694 3591 2746
rect 3591 2694 3621 2746
rect 3645 2694 3655 2746
rect 3655 2694 3701 2746
rect 3405 2692 3461 2694
rect 3485 2692 3541 2694
rect 3565 2692 3621 2694
rect 3645 2692 3701 2694
rect 1490 2216 1546 2272
rect 5854 20698 5910 20700
rect 5934 20698 5990 20700
rect 6014 20698 6070 20700
rect 6094 20698 6150 20700
rect 5854 20646 5900 20698
rect 5900 20646 5910 20698
rect 5934 20646 5964 20698
rect 5964 20646 5976 20698
rect 5976 20646 5990 20698
rect 6014 20646 6028 20698
rect 6028 20646 6040 20698
rect 6040 20646 6070 20698
rect 6094 20646 6104 20698
rect 6104 20646 6150 20698
rect 5854 20644 5910 20646
rect 5934 20644 5990 20646
rect 6014 20644 6070 20646
rect 6094 20644 6150 20646
rect 5854 19610 5910 19612
rect 5934 19610 5990 19612
rect 6014 19610 6070 19612
rect 6094 19610 6150 19612
rect 5854 19558 5900 19610
rect 5900 19558 5910 19610
rect 5934 19558 5964 19610
rect 5964 19558 5976 19610
rect 5976 19558 5990 19610
rect 6014 19558 6028 19610
rect 6028 19558 6040 19610
rect 6040 19558 6070 19610
rect 6094 19558 6104 19610
rect 6104 19558 6150 19610
rect 5854 19556 5910 19558
rect 5934 19556 5990 19558
rect 6014 19556 6070 19558
rect 6094 19556 6150 19558
rect 5854 18522 5910 18524
rect 5934 18522 5990 18524
rect 6014 18522 6070 18524
rect 6094 18522 6150 18524
rect 5854 18470 5900 18522
rect 5900 18470 5910 18522
rect 5934 18470 5964 18522
rect 5964 18470 5976 18522
rect 5976 18470 5990 18522
rect 6014 18470 6028 18522
rect 6028 18470 6040 18522
rect 6040 18470 6070 18522
rect 6094 18470 6104 18522
rect 6104 18470 6150 18522
rect 5854 18468 5910 18470
rect 5934 18468 5990 18470
rect 6014 18468 6070 18470
rect 6094 18468 6150 18470
rect 5854 17434 5910 17436
rect 5934 17434 5990 17436
rect 6014 17434 6070 17436
rect 6094 17434 6150 17436
rect 5854 17382 5900 17434
rect 5900 17382 5910 17434
rect 5934 17382 5964 17434
rect 5964 17382 5976 17434
rect 5976 17382 5990 17434
rect 6014 17382 6028 17434
rect 6028 17382 6040 17434
rect 6040 17382 6070 17434
rect 6094 17382 6104 17434
rect 6104 17382 6150 17434
rect 5854 17380 5910 17382
rect 5934 17380 5990 17382
rect 6014 17380 6070 17382
rect 6094 17380 6150 17382
rect 5854 16346 5910 16348
rect 5934 16346 5990 16348
rect 6014 16346 6070 16348
rect 6094 16346 6150 16348
rect 5854 16294 5900 16346
rect 5900 16294 5910 16346
rect 5934 16294 5964 16346
rect 5964 16294 5976 16346
rect 5976 16294 5990 16346
rect 6014 16294 6028 16346
rect 6028 16294 6040 16346
rect 6040 16294 6070 16346
rect 6094 16294 6104 16346
rect 6104 16294 6150 16346
rect 5854 16292 5910 16294
rect 5934 16292 5990 16294
rect 6014 16292 6070 16294
rect 6094 16292 6150 16294
rect 5854 15258 5910 15260
rect 5934 15258 5990 15260
rect 6014 15258 6070 15260
rect 6094 15258 6150 15260
rect 5854 15206 5900 15258
rect 5900 15206 5910 15258
rect 5934 15206 5964 15258
rect 5964 15206 5976 15258
rect 5976 15206 5990 15258
rect 6014 15206 6028 15258
rect 6028 15206 6040 15258
rect 6040 15206 6070 15258
rect 6094 15206 6104 15258
rect 6104 15206 6150 15258
rect 5854 15204 5910 15206
rect 5934 15204 5990 15206
rect 6014 15204 6070 15206
rect 6094 15204 6150 15206
rect 5854 14170 5910 14172
rect 5934 14170 5990 14172
rect 6014 14170 6070 14172
rect 6094 14170 6150 14172
rect 5854 14118 5900 14170
rect 5900 14118 5910 14170
rect 5934 14118 5964 14170
rect 5964 14118 5976 14170
rect 5976 14118 5990 14170
rect 6014 14118 6028 14170
rect 6028 14118 6040 14170
rect 6040 14118 6070 14170
rect 6094 14118 6104 14170
rect 6104 14118 6150 14170
rect 5854 14116 5910 14118
rect 5934 14116 5990 14118
rect 6014 14116 6070 14118
rect 6094 14116 6150 14118
rect 5854 13082 5910 13084
rect 5934 13082 5990 13084
rect 6014 13082 6070 13084
rect 6094 13082 6150 13084
rect 5854 13030 5900 13082
rect 5900 13030 5910 13082
rect 5934 13030 5964 13082
rect 5964 13030 5976 13082
rect 5976 13030 5990 13082
rect 6014 13030 6028 13082
rect 6028 13030 6040 13082
rect 6040 13030 6070 13082
rect 6094 13030 6104 13082
rect 6104 13030 6150 13082
rect 5854 13028 5910 13030
rect 5934 13028 5990 13030
rect 6014 13028 6070 13030
rect 6094 13028 6150 13030
rect 5854 11994 5910 11996
rect 5934 11994 5990 11996
rect 6014 11994 6070 11996
rect 6094 11994 6150 11996
rect 5854 11942 5900 11994
rect 5900 11942 5910 11994
rect 5934 11942 5964 11994
rect 5964 11942 5976 11994
rect 5976 11942 5990 11994
rect 6014 11942 6028 11994
rect 6028 11942 6040 11994
rect 6040 11942 6070 11994
rect 6094 11942 6104 11994
rect 6104 11942 6150 11994
rect 5854 11940 5910 11942
rect 5934 11940 5990 11942
rect 6014 11940 6070 11942
rect 6094 11940 6150 11942
rect 5854 10906 5910 10908
rect 5934 10906 5990 10908
rect 6014 10906 6070 10908
rect 6094 10906 6150 10908
rect 5854 10854 5900 10906
rect 5900 10854 5910 10906
rect 5934 10854 5964 10906
rect 5964 10854 5976 10906
rect 5976 10854 5990 10906
rect 6014 10854 6028 10906
rect 6028 10854 6040 10906
rect 6040 10854 6070 10906
rect 6094 10854 6104 10906
rect 6104 10854 6150 10906
rect 5854 10852 5910 10854
rect 5934 10852 5990 10854
rect 6014 10852 6070 10854
rect 6094 10852 6150 10854
rect 5854 9818 5910 9820
rect 5934 9818 5990 9820
rect 6014 9818 6070 9820
rect 6094 9818 6150 9820
rect 5854 9766 5900 9818
rect 5900 9766 5910 9818
rect 5934 9766 5964 9818
rect 5964 9766 5976 9818
rect 5976 9766 5990 9818
rect 6014 9766 6028 9818
rect 6028 9766 6040 9818
rect 6040 9766 6070 9818
rect 6094 9766 6104 9818
rect 6104 9766 6150 9818
rect 5854 9764 5910 9766
rect 5934 9764 5990 9766
rect 6014 9764 6070 9766
rect 6094 9764 6150 9766
rect 4894 6160 4950 6216
rect 5854 8730 5910 8732
rect 5934 8730 5990 8732
rect 6014 8730 6070 8732
rect 6094 8730 6150 8732
rect 5854 8678 5900 8730
rect 5900 8678 5910 8730
rect 5934 8678 5964 8730
rect 5964 8678 5976 8730
rect 5976 8678 5990 8730
rect 6014 8678 6028 8730
rect 6028 8678 6040 8730
rect 6040 8678 6070 8730
rect 6094 8678 6104 8730
rect 6104 8678 6150 8730
rect 5854 8676 5910 8678
rect 5934 8676 5990 8678
rect 6014 8676 6070 8678
rect 6094 8676 6150 8678
rect 8304 21242 8360 21244
rect 8384 21242 8440 21244
rect 8464 21242 8520 21244
rect 8544 21242 8600 21244
rect 8304 21190 8350 21242
rect 8350 21190 8360 21242
rect 8384 21190 8414 21242
rect 8414 21190 8426 21242
rect 8426 21190 8440 21242
rect 8464 21190 8478 21242
rect 8478 21190 8490 21242
rect 8490 21190 8520 21242
rect 8544 21190 8554 21242
rect 8554 21190 8600 21242
rect 8304 21188 8360 21190
rect 8384 21188 8440 21190
rect 8464 21188 8520 21190
rect 8544 21188 8600 21190
rect 8304 20154 8360 20156
rect 8384 20154 8440 20156
rect 8464 20154 8520 20156
rect 8544 20154 8600 20156
rect 8304 20102 8350 20154
rect 8350 20102 8360 20154
rect 8384 20102 8414 20154
rect 8414 20102 8426 20154
rect 8426 20102 8440 20154
rect 8464 20102 8478 20154
rect 8478 20102 8490 20154
rect 8490 20102 8520 20154
rect 8544 20102 8554 20154
rect 8554 20102 8600 20154
rect 8304 20100 8360 20102
rect 8384 20100 8440 20102
rect 8464 20100 8520 20102
rect 8544 20100 8600 20102
rect 8304 19066 8360 19068
rect 8384 19066 8440 19068
rect 8464 19066 8520 19068
rect 8544 19066 8600 19068
rect 8304 19014 8350 19066
rect 8350 19014 8360 19066
rect 8384 19014 8414 19066
rect 8414 19014 8426 19066
rect 8426 19014 8440 19066
rect 8464 19014 8478 19066
rect 8478 19014 8490 19066
rect 8490 19014 8520 19066
rect 8544 19014 8554 19066
rect 8554 19014 8600 19066
rect 8304 19012 8360 19014
rect 8384 19012 8440 19014
rect 8464 19012 8520 19014
rect 8544 19012 8600 19014
rect 8304 17978 8360 17980
rect 8384 17978 8440 17980
rect 8464 17978 8520 17980
rect 8544 17978 8600 17980
rect 8304 17926 8350 17978
rect 8350 17926 8360 17978
rect 8384 17926 8414 17978
rect 8414 17926 8426 17978
rect 8426 17926 8440 17978
rect 8464 17926 8478 17978
rect 8478 17926 8490 17978
rect 8490 17926 8520 17978
rect 8544 17926 8554 17978
rect 8554 17926 8600 17978
rect 8304 17924 8360 17926
rect 8384 17924 8440 17926
rect 8464 17924 8520 17926
rect 8544 17924 8600 17926
rect 8304 16890 8360 16892
rect 8384 16890 8440 16892
rect 8464 16890 8520 16892
rect 8544 16890 8600 16892
rect 8304 16838 8350 16890
rect 8350 16838 8360 16890
rect 8384 16838 8414 16890
rect 8414 16838 8426 16890
rect 8426 16838 8440 16890
rect 8464 16838 8478 16890
rect 8478 16838 8490 16890
rect 8490 16838 8520 16890
rect 8544 16838 8554 16890
rect 8554 16838 8600 16890
rect 8304 16836 8360 16838
rect 8384 16836 8440 16838
rect 8464 16836 8520 16838
rect 8544 16836 8600 16838
rect 8304 15802 8360 15804
rect 8384 15802 8440 15804
rect 8464 15802 8520 15804
rect 8544 15802 8600 15804
rect 8304 15750 8350 15802
rect 8350 15750 8360 15802
rect 8384 15750 8414 15802
rect 8414 15750 8426 15802
rect 8426 15750 8440 15802
rect 8464 15750 8478 15802
rect 8478 15750 8490 15802
rect 8490 15750 8520 15802
rect 8544 15750 8554 15802
rect 8554 15750 8600 15802
rect 8304 15748 8360 15750
rect 8384 15748 8440 15750
rect 8464 15748 8520 15750
rect 8544 15748 8600 15750
rect 8304 14714 8360 14716
rect 8384 14714 8440 14716
rect 8464 14714 8520 14716
rect 8544 14714 8600 14716
rect 8304 14662 8350 14714
rect 8350 14662 8360 14714
rect 8384 14662 8414 14714
rect 8414 14662 8426 14714
rect 8426 14662 8440 14714
rect 8464 14662 8478 14714
rect 8478 14662 8490 14714
rect 8490 14662 8520 14714
rect 8544 14662 8554 14714
rect 8554 14662 8600 14714
rect 8304 14660 8360 14662
rect 8384 14660 8440 14662
rect 8464 14660 8520 14662
rect 8544 14660 8600 14662
rect 8304 13626 8360 13628
rect 8384 13626 8440 13628
rect 8464 13626 8520 13628
rect 8544 13626 8600 13628
rect 8304 13574 8350 13626
rect 8350 13574 8360 13626
rect 8384 13574 8414 13626
rect 8414 13574 8426 13626
rect 8426 13574 8440 13626
rect 8464 13574 8478 13626
rect 8478 13574 8490 13626
rect 8490 13574 8520 13626
rect 8544 13574 8554 13626
rect 8554 13574 8600 13626
rect 8304 13572 8360 13574
rect 8384 13572 8440 13574
rect 8464 13572 8520 13574
rect 8544 13572 8600 13574
rect 8304 12538 8360 12540
rect 8384 12538 8440 12540
rect 8464 12538 8520 12540
rect 8544 12538 8600 12540
rect 8304 12486 8350 12538
rect 8350 12486 8360 12538
rect 8384 12486 8414 12538
rect 8414 12486 8426 12538
rect 8426 12486 8440 12538
rect 8464 12486 8478 12538
rect 8478 12486 8490 12538
rect 8490 12486 8520 12538
rect 8544 12486 8554 12538
rect 8554 12486 8600 12538
rect 8304 12484 8360 12486
rect 8384 12484 8440 12486
rect 8464 12484 8520 12486
rect 8544 12484 8600 12486
rect 8304 11450 8360 11452
rect 8384 11450 8440 11452
rect 8464 11450 8520 11452
rect 8544 11450 8600 11452
rect 8304 11398 8350 11450
rect 8350 11398 8360 11450
rect 8384 11398 8414 11450
rect 8414 11398 8426 11450
rect 8426 11398 8440 11450
rect 8464 11398 8478 11450
rect 8478 11398 8490 11450
rect 8490 11398 8520 11450
rect 8544 11398 8554 11450
rect 8554 11398 8600 11450
rect 8304 11396 8360 11398
rect 8384 11396 8440 11398
rect 8464 11396 8520 11398
rect 8544 11396 8600 11398
rect 5854 7642 5910 7644
rect 5934 7642 5990 7644
rect 6014 7642 6070 7644
rect 6094 7642 6150 7644
rect 5854 7590 5900 7642
rect 5900 7590 5910 7642
rect 5934 7590 5964 7642
rect 5964 7590 5976 7642
rect 5976 7590 5990 7642
rect 6014 7590 6028 7642
rect 6028 7590 6040 7642
rect 6040 7590 6070 7642
rect 6094 7590 6104 7642
rect 6104 7590 6150 7642
rect 5854 7588 5910 7590
rect 5934 7588 5990 7590
rect 6014 7588 6070 7590
rect 6094 7588 6150 7590
rect 5854 6554 5910 6556
rect 5934 6554 5990 6556
rect 6014 6554 6070 6556
rect 6094 6554 6150 6556
rect 5854 6502 5900 6554
rect 5900 6502 5910 6554
rect 5934 6502 5964 6554
rect 5964 6502 5976 6554
rect 5976 6502 5990 6554
rect 6014 6502 6028 6554
rect 6028 6502 6040 6554
rect 6040 6502 6070 6554
rect 6094 6502 6104 6554
rect 6104 6502 6150 6554
rect 5854 6500 5910 6502
rect 5934 6500 5990 6502
rect 6014 6500 6070 6502
rect 6094 6500 6150 6502
rect 5854 5466 5910 5468
rect 5934 5466 5990 5468
rect 6014 5466 6070 5468
rect 6094 5466 6150 5468
rect 5854 5414 5900 5466
rect 5900 5414 5910 5466
rect 5934 5414 5964 5466
rect 5964 5414 5976 5466
rect 5976 5414 5990 5466
rect 6014 5414 6028 5466
rect 6028 5414 6040 5466
rect 6040 5414 6070 5466
rect 6094 5414 6104 5466
rect 6104 5414 6150 5466
rect 5854 5412 5910 5414
rect 5934 5412 5990 5414
rect 6014 5412 6070 5414
rect 6094 5412 6150 5414
rect 5854 4378 5910 4380
rect 5934 4378 5990 4380
rect 6014 4378 6070 4380
rect 6094 4378 6150 4380
rect 5854 4326 5900 4378
rect 5900 4326 5910 4378
rect 5934 4326 5964 4378
rect 5964 4326 5976 4378
rect 5976 4326 5990 4378
rect 6014 4326 6028 4378
rect 6028 4326 6040 4378
rect 6040 4326 6070 4378
rect 6094 4326 6104 4378
rect 6104 4326 6150 4378
rect 5854 4324 5910 4326
rect 5934 4324 5990 4326
rect 6014 4324 6070 4326
rect 6094 4324 6150 4326
rect 5854 3290 5910 3292
rect 5934 3290 5990 3292
rect 6014 3290 6070 3292
rect 6094 3290 6150 3292
rect 5854 3238 5900 3290
rect 5900 3238 5910 3290
rect 5934 3238 5964 3290
rect 5964 3238 5976 3290
rect 5976 3238 5990 3290
rect 6014 3238 6028 3290
rect 6028 3238 6040 3290
rect 6040 3238 6070 3290
rect 6094 3238 6104 3290
rect 6104 3238 6150 3290
rect 5854 3236 5910 3238
rect 5934 3236 5990 3238
rect 6014 3236 6070 3238
rect 6094 3236 6150 3238
rect 8304 10362 8360 10364
rect 8384 10362 8440 10364
rect 8464 10362 8520 10364
rect 8544 10362 8600 10364
rect 8304 10310 8350 10362
rect 8350 10310 8360 10362
rect 8384 10310 8414 10362
rect 8414 10310 8426 10362
rect 8426 10310 8440 10362
rect 8464 10310 8478 10362
rect 8478 10310 8490 10362
rect 8490 10310 8520 10362
rect 8544 10310 8554 10362
rect 8554 10310 8600 10362
rect 8304 10308 8360 10310
rect 8384 10308 8440 10310
rect 8464 10308 8520 10310
rect 8544 10308 8600 10310
rect 8304 9274 8360 9276
rect 8384 9274 8440 9276
rect 8464 9274 8520 9276
rect 8544 9274 8600 9276
rect 8304 9222 8350 9274
rect 8350 9222 8360 9274
rect 8384 9222 8414 9274
rect 8414 9222 8426 9274
rect 8426 9222 8440 9274
rect 8464 9222 8478 9274
rect 8478 9222 8490 9274
rect 8490 9222 8520 9274
rect 8544 9222 8554 9274
rect 8554 9222 8600 9274
rect 8304 9220 8360 9222
rect 8384 9220 8440 9222
rect 8464 9220 8520 9222
rect 8544 9220 8600 9222
rect 8304 8186 8360 8188
rect 8384 8186 8440 8188
rect 8464 8186 8520 8188
rect 8544 8186 8600 8188
rect 8304 8134 8350 8186
rect 8350 8134 8360 8186
rect 8384 8134 8414 8186
rect 8414 8134 8426 8186
rect 8426 8134 8440 8186
rect 8464 8134 8478 8186
rect 8478 8134 8490 8186
rect 8490 8134 8520 8186
rect 8544 8134 8554 8186
rect 8554 8134 8600 8186
rect 8304 8132 8360 8134
rect 8384 8132 8440 8134
rect 8464 8132 8520 8134
rect 8544 8132 8600 8134
rect 8304 7098 8360 7100
rect 8384 7098 8440 7100
rect 8464 7098 8520 7100
rect 8544 7098 8600 7100
rect 8304 7046 8350 7098
rect 8350 7046 8360 7098
rect 8384 7046 8414 7098
rect 8414 7046 8426 7098
rect 8426 7046 8440 7098
rect 8464 7046 8478 7098
rect 8478 7046 8490 7098
rect 8490 7046 8520 7098
rect 8544 7046 8554 7098
rect 8554 7046 8600 7098
rect 8304 7044 8360 7046
rect 8384 7044 8440 7046
rect 8464 7044 8520 7046
rect 8544 7044 8600 7046
rect 8304 6010 8360 6012
rect 8384 6010 8440 6012
rect 8464 6010 8520 6012
rect 8544 6010 8600 6012
rect 8304 5958 8350 6010
rect 8350 5958 8360 6010
rect 8384 5958 8414 6010
rect 8414 5958 8426 6010
rect 8426 5958 8440 6010
rect 8464 5958 8478 6010
rect 8478 5958 8490 6010
rect 8490 5958 8520 6010
rect 8544 5958 8554 6010
rect 8554 5958 8600 6010
rect 8304 5956 8360 5958
rect 8384 5956 8440 5958
rect 8464 5956 8520 5958
rect 8544 5956 8600 5958
rect 8304 4922 8360 4924
rect 8384 4922 8440 4924
rect 8464 4922 8520 4924
rect 8544 4922 8600 4924
rect 8304 4870 8350 4922
rect 8350 4870 8360 4922
rect 8384 4870 8414 4922
rect 8414 4870 8426 4922
rect 8426 4870 8440 4922
rect 8464 4870 8478 4922
rect 8478 4870 8490 4922
rect 8490 4870 8520 4922
rect 8544 4870 8554 4922
rect 8554 4870 8600 4922
rect 8304 4868 8360 4870
rect 8384 4868 8440 4870
rect 8464 4868 8520 4870
rect 8544 4868 8600 4870
rect 8304 3834 8360 3836
rect 8384 3834 8440 3836
rect 8464 3834 8520 3836
rect 8544 3834 8600 3836
rect 8304 3782 8350 3834
rect 8350 3782 8360 3834
rect 8384 3782 8414 3834
rect 8414 3782 8426 3834
rect 8426 3782 8440 3834
rect 8464 3782 8478 3834
rect 8478 3782 8490 3834
rect 8490 3782 8520 3834
rect 8544 3782 8554 3834
rect 8554 3782 8600 3834
rect 8304 3780 8360 3782
rect 8384 3780 8440 3782
rect 8464 3780 8520 3782
rect 8544 3780 8600 3782
rect 8304 2746 8360 2748
rect 8384 2746 8440 2748
rect 8464 2746 8520 2748
rect 8544 2746 8600 2748
rect 8304 2694 8350 2746
rect 8350 2694 8360 2746
rect 8384 2694 8414 2746
rect 8414 2694 8426 2746
rect 8426 2694 8440 2746
rect 8464 2694 8478 2746
rect 8478 2694 8490 2746
rect 8490 2694 8520 2746
rect 8544 2694 8554 2746
rect 8554 2694 8600 2746
rect 8304 2692 8360 2694
rect 8384 2692 8440 2694
rect 8464 2692 8520 2694
rect 8544 2692 8600 2694
rect 10753 20698 10809 20700
rect 10833 20698 10889 20700
rect 10913 20698 10969 20700
rect 10993 20698 11049 20700
rect 10753 20646 10799 20698
rect 10799 20646 10809 20698
rect 10833 20646 10863 20698
rect 10863 20646 10875 20698
rect 10875 20646 10889 20698
rect 10913 20646 10927 20698
rect 10927 20646 10939 20698
rect 10939 20646 10969 20698
rect 10993 20646 11003 20698
rect 11003 20646 11049 20698
rect 10753 20644 10809 20646
rect 10833 20644 10889 20646
rect 10913 20644 10969 20646
rect 10993 20644 11049 20646
rect 13203 21242 13259 21244
rect 13283 21242 13339 21244
rect 13363 21242 13419 21244
rect 13443 21242 13499 21244
rect 13203 21190 13249 21242
rect 13249 21190 13259 21242
rect 13283 21190 13313 21242
rect 13313 21190 13325 21242
rect 13325 21190 13339 21242
rect 13363 21190 13377 21242
rect 13377 21190 13389 21242
rect 13389 21190 13419 21242
rect 13443 21190 13453 21242
rect 13453 21190 13499 21242
rect 13203 21188 13259 21190
rect 13283 21188 13339 21190
rect 13363 21188 13419 21190
rect 13443 21188 13499 21190
rect 10753 19610 10809 19612
rect 10833 19610 10889 19612
rect 10913 19610 10969 19612
rect 10993 19610 11049 19612
rect 10753 19558 10799 19610
rect 10799 19558 10809 19610
rect 10833 19558 10863 19610
rect 10863 19558 10875 19610
rect 10875 19558 10889 19610
rect 10913 19558 10927 19610
rect 10927 19558 10939 19610
rect 10939 19558 10969 19610
rect 10993 19558 11003 19610
rect 11003 19558 11049 19610
rect 10753 19556 10809 19558
rect 10833 19556 10889 19558
rect 10913 19556 10969 19558
rect 10993 19556 11049 19558
rect 10753 18522 10809 18524
rect 10833 18522 10889 18524
rect 10913 18522 10969 18524
rect 10993 18522 11049 18524
rect 10753 18470 10799 18522
rect 10799 18470 10809 18522
rect 10833 18470 10863 18522
rect 10863 18470 10875 18522
rect 10875 18470 10889 18522
rect 10913 18470 10927 18522
rect 10927 18470 10939 18522
rect 10939 18470 10969 18522
rect 10993 18470 11003 18522
rect 11003 18470 11049 18522
rect 10753 18468 10809 18470
rect 10833 18468 10889 18470
rect 10913 18468 10969 18470
rect 10993 18468 11049 18470
rect 13203 20154 13259 20156
rect 13283 20154 13339 20156
rect 13363 20154 13419 20156
rect 13443 20154 13499 20156
rect 13203 20102 13249 20154
rect 13249 20102 13259 20154
rect 13283 20102 13313 20154
rect 13313 20102 13325 20154
rect 13325 20102 13339 20154
rect 13363 20102 13377 20154
rect 13377 20102 13389 20154
rect 13389 20102 13419 20154
rect 13443 20102 13453 20154
rect 13453 20102 13499 20154
rect 13203 20100 13259 20102
rect 13283 20100 13339 20102
rect 13363 20100 13419 20102
rect 13443 20100 13499 20102
rect 13203 19066 13259 19068
rect 13283 19066 13339 19068
rect 13363 19066 13419 19068
rect 13443 19066 13499 19068
rect 13203 19014 13249 19066
rect 13249 19014 13259 19066
rect 13283 19014 13313 19066
rect 13313 19014 13325 19066
rect 13325 19014 13339 19066
rect 13363 19014 13377 19066
rect 13377 19014 13389 19066
rect 13389 19014 13419 19066
rect 13443 19014 13453 19066
rect 13453 19014 13499 19066
rect 13203 19012 13259 19014
rect 13283 19012 13339 19014
rect 13363 19012 13419 19014
rect 13443 19012 13499 19014
rect 10753 17434 10809 17436
rect 10833 17434 10889 17436
rect 10913 17434 10969 17436
rect 10993 17434 11049 17436
rect 10753 17382 10799 17434
rect 10799 17382 10809 17434
rect 10833 17382 10863 17434
rect 10863 17382 10875 17434
rect 10875 17382 10889 17434
rect 10913 17382 10927 17434
rect 10927 17382 10939 17434
rect 10939 17382 10969 17434
rect 10993 17382 11003 17434
rect 11003 17382 11049 17434
rect 10753 17380 10809 17382
rect 10833 17380 10889 17382
rect 10913 17380 10969 17382
rect 10993 17380 11049 17382
rect 10753 16346 10809 16348
rect 10833 16346 10889 16348
rect 10913 16346 10969 16348
rect 10993 16346 11049 16348
rect 10753 16294 10799 16346
rect 10799 16294 10809 16346
rect 10833 16294 10863 16346
rect 10863 16294 10875 16346
rect 10875 16294 10889 16346
rect 10913 16294 10927 16346
rect 10927 16294 10939 16346
rect 10939 16294 10969 16346
rect 10993 16294 11003 16346
rect 11003 16294 11049 16346
rect 10753 16292 10809 16294
rect 10833 16292 10889 16294
rect 10913 16292 10969 16294
rect 10993 16292 11049 16294
rect 10753 15258 10809 15260
rect 10833 15258 10889 15260
rect 10913 15258 10969 15260
rect 10993 15258 11049 15260
rect 10753 15206 10799 15258
rect 10799 15206 10809 15258
rect 10833 15206 10863 15258
rect 10863 15206 10875 15258
rect 10875 15206 10889 15258
rect 10913 15206 10927 15258
rect 10927 15206 10939 15258
rect 10939 15206 10969 15258
rect 10993 15206 11003 15258
rect 11003 15206 11049 15258
rect 10753 15204 10809 15206
rect 10833 15204 10889 15206
rect 10913 15204 10969 15206
rect 10993 15204 11049 15206
rect 10753 14170 10809 14172
rect 10833 14170 10889 14172
rect 10913 14170 10969 14172
rect 10993 14170 11049 14172
rect 10753 14118 10799 14170
rect 10799 14118 10809 14170
rect 10833 14118 10863 14170
rect 10863 14118 10875 14170
rect 10875 14118 10889 14170
rect 10913 14118 10927 14170
rect 10927 14118 10939 14170
rect 10939 14118 10969 14170
rect 10993 14118 11003 14170
rect 11003 14118 11049 14170
rect 10753 14116 10809 14118
rect 10833 14116 10889 14118
rect 10913 14116 10969 14118
rect 10993 14116 11049 14118
rect 10753 13082 10809 13084
rect 10833 13082 10889 13084
rect 10913 13082 10969 13084
rect 10993 13082 11049 13084
rect 10753 13030 10799 13082
rect 10799 13030 10809 13082
rect 10833 13030 10863 13082
rect 10863 13030 10875 13082
rect 10875 13030 10889 13082
rect 10913 13030 10927 13082
rect 10927 13030 10939 13082
rect 10939 13030 10969 13082
rect 10993 13030 11003 13082
rect 11003 13030 11049 13082
rect 10753 13028 10809 13030
rect 10833 13028 10889 13030
rect 10913 13028 10969 13030
rect 10993 13028 11049 13030
rect 13203 17978 13259 17980
rect 13283 17978 13339 17980
rect 13363 17978 13419 17980
rect 13443 17978 13499 17980
rect 13203 17926 13249 17978
rect 13249 17926 13259 17978
rect 13283 17926 13313 17978
rect 13313 17926 13325 17978
rect 13325 17926 13339 17978
rect 13363 17926 13377 17978
rect 13377 17926 13389 17978
rect 13389 17926 13419 17978
rect 13443 17926 13453 17978
rect 13453 17926 13499 17978
rect 13203 17924 13259 17926
rect 13283 17924 13339 17926
rect 13363 17924 13419 17926
rect 13443 17924 13499 17926
rect 13203 16890 13259 16892
rect 13283 16890 13339 16892
rect 13363 16890 13419 16892
rect 13443 16890 13499 16892
rect 13203 16838 13249 16890
rect 13249 16838 13259 16890
rect 13283 16838 13313 16890
rect 13313 16838 13325 16890
rect 13325 16838 13339 16890
rect 13363 16838 13377 16890
rect 13377 16838 13389 16890
rect 13389 16838 13419 16890
rect 13443 16838 13453 16890
rect 13453 16838 13499 16890
rect 13203 16836 13259 16838
rect 13283 16836 13339 16838
rect 13363 16836 13419 16838
rect 13443 16836 13499 16838
rect 13203 15802 13259 15804
rect 13283 15802 13339 15804
rect 13363 15802 13419 15804
rect 13443 15802 13499 15804
rect 13203 15750 13249 15802
rect 13249 15750 13259 15802
rect 13283 15750 13313 15802
rect 13313 15750 13325 15802
rect 13325 15750 13339 15802
rect 13363 15750 13377 15802
rect 13377 15750 13389 15802
rect 13389 15750 13419 15802
rect 13443 15750 13453 15802
rect 13453 15750 13499 15802
rect 13203 15748 13259 15750
rect 13283 15748 13339 15750
rect 13363 15748 13419 15750
rect 13443 15748 13499 15750
rect 13203 14714 13259 14716
rect 13283 14714 13339 14716
rect 13363 14714 13419 14716
rect 13443 14714 13499 14716
rect 13203 14662 13249 14714
rect 13249 14662 13259 14714
rect 13283 14662 13313 14714
rect 13313 14662 13325 14714
rect 13325 14662 13339 14714
rect 13363 14662 13377 14714
rect 13377 14662 13389 14714
rect 13389 14662 13419 14714
rect 13443 14662 13453 14714
rect 13453 14662 13499 14714
rect 13203 14660 13259 14662
rect 13283 14660 13339 14662
rect 13363 14660 13419 14662
rect 13443 14660 13499 14662
rect 13203 13626 13259 13628
rect 13283 13626 13339 13628
rect 13363 13626 13419 13628
rect 13443 13626 13499 13628
rect 13203 13574 13249 13626
rect 13249 13574 13259 13626
rect 13283 13574 13313 13626
rect 13313 13574 13325 13626
rect 13325 13574 13339 13626
rect 13363 13574 13377 13626
rect 13377 13574 13389 13626
rect 13389 13574 13419 13626
rect 13443 13574 13453 13626
rect 13453 13574 13499 13626
rect 13203 13572 13259 13574
rect 13283 13572 13339 13574
rect 13363 13572 13419 13574
rect 13443 13572 13499 13574
rect 13203 12538 13259 12540
rect 13283 12538 13339 12540
rect 13363 12538 13419 12540
rect 13443 12538 13499 12540
rect 13203 12486 13249 12538
rect 13249 12486 13259 12538
rect 13283 12486 13313 12538
rect 13313 12486 13325 12538
rect 13325 12486 13339 12538
rect 13363 12486 13377 12538
rect 13377 12486 13389 12538
rect 13389 12486 13419 12538
rect 13443 12486 13453 12538
rect 13453 12486 13499 12538
rect 13203 12484 13259 12486
rect 13283 12484 13339 12486
rect 13363 12484 13419 12486
rect 13443 12484 13499 12486
rect 10753 11994 10809 11996
rect 10833 11994 10889 11996
rect 10913 11994 10969 11996
rect 10993 11994 11049 11996
rect 10753 11942 10799 11994
rect 10799 11942 10809 11994
rect 10833 11942 10863 11994
rect 10863 11942 10875 11994
rect 10875 11942 10889 11994
rect 10913 11942 10927 11994
rect 10927 11942 10939 11994
rect 10939 11942 10969 11994
rect 10993 11942 11003 11994
rect 11003 11942 11049 11994
rect 10753 11940 10809 11942
rect 10833 11940 10889 11942
rect 10913 11940 10969 11942
rect 10993 11940 11049 11942
rect 10753 10906 10809 10908
rect 10833 10906 10889 10908
rect 10913 10906 10969 10908
rect 10993 10906 11049 10908
rect 10753 10854 10799 10906
rect 10799 10854 10809 10906
rect 10833 10854 10863 10906
rect 10863 10854 10875 10906
rect 10875 10854 10889 10906
rect 10913 10854 10927 10906
rect 10927 10854 10939 10906
rect 10939 10854 10969 10906
rect 10993 10854 11003 10906
rect 11003 10854 11049 10906
rect 10753 10852 10809 10854
rect 10833 10852 10889 10854
rect 10913 10852 10969 10854
rect 10993 10852 11049 10854
rect 10753 9818 10809 9820
rect 10833 9818 10889 9820
rect 10913 9818 10969 9820
rect 10993 9818 11049 9820
rect 10753 9766 10799 9818
rect 10799 9766 10809 9818
rect 10833 9766 10863 9818
rect 10863 9766 10875 9818
rect 10875 9766 10889 9818
rect 10913 9766 10927 9818
rect 10927 9766 10939 9818
rect 10939 9766 10969 9818
rect 10993 9766 11003 9818
rect 11003 9766 11049 9818
rect 10753 9764 10809 9766
rect 10833 9764 10889 9766
rect 10913 9764 10969 9766
rect 10993 9764 11049 9766
rect 10753 8730 10809 8732
rect 10833 8730 10889 8732
rect 10913 8730 10969 8732
rect 10993 8730 11049 8732
rect 10753 8678 10799 8730
rect 10799 8678 10809 8730
rect 10833 8678 10863 8730
rect 10863 8678 10875 8730
rect 10875 8678 10889 8730
rect 10913 8678 10927 8730
rect 10927 8678 10939 8730
rect 10939 8678 10969 8730
rect 10993 8678 11003 8730
rect 11003 8678 11049 8730
rect 10753 8676 10809 8678
rect 10833 8676 10889 8678
rect 10913 8676 10969 8678
rect 10993 8676 11049 8678
rect 10753 7642 10809 7644
rect 10833 7642 10889 7644
rect 10913 7642 10969 7644
rect 10993 7642 11049 7644
rect 10753 7590 10799 7642
rect 10799 7590 10809 7642
rect 10833 7590 10863 7642
rect 10863 7590 10875 7642
rect 10875 7590 10889 7642
rect 10913 7590 10927 7642
rect 10927 7590 10939 7642
rect 10939 7590 10969 7642
rect 10993 7590 11003 7642
rect 11003 7590 11049 7642
rect 10753 7588 10809 7590
rect 10833 7588 10889 7590
rect 10913 7588 10969 7590
rect 10993 7588 11049 7590
rect 13203 11450 13259 11452
rect 13283 11450 13339 11452
rect 13363 11450 13419 11452
rect 13443 11450 13499 11452
rect 13203 11398 13249 11450
rect 13249 11398 13259 11450
rect 13283 11398 13313 11450
rect 13313 11398 13325 11450
rect 13325 11398 13339 11450
rect 13363 11398 13377 11450
rect 13377 11398 13389 11450
rect 13389 11398 13419 11450
rect 13443 11398 13453 11450
rect 13453 11398 13499 11450
rect 13203 11396 13259 11398
rect 13283 11396 13339 11398
rect 13363 11396 13419 11398
rect 13443 11396 13499 11398
rect 13203 10362 13259 10364
rect 13283 10362 13339 10364
rect 13363 10362 13419 10364
rect 13443 10362 13499 10364
rect 13203 10310 13249 10362
rect 13249 10310 13259 10362
rect 13283 10310 13313 10362
rect 13313 10310 13325 10362
rect 13325 10310 13339 10362
rect 13363 10310 13377 10362
rect 13377 10310 13389 10362
rect 13389 10310 13419 10362
rect 13443 10310 13453 10362
rect 13453 10310 13499 10362
rect 13203 10308 13259 10310
rect 13283 10308 13339 10310
rect 13363 10308 13419 10310
rect 13443 10308 13499 10310
rect 13203 9274 13259 9276
rect 13283 9274 13339 9276
rect 13363 9274 13419 9276
rect 13443 9274 13499 9276
rect 13203 9222 13249 9274
rect 13249 9222 13259 9274
rect 13283 9222 13313 9274
rect 13313 9222 13325 9274
rect 13325 9222 13339 9274
rect 13363 9222 13377 9274
rect 13377 9222 13389 9274
rect 13389 9222 13419 9274
rect 13443 9222 13453 9274
rect 13453 9222 13499 9274
rect 13203 9220 13259 9222
rect 13283 9220 13339 9222
rect 13363 9220 13419 9222
rect 13443 9220 13499 9222
rect 13203 8186 13259 8188
rect 13283 8186 13339 8188
rect 13363 8186 13419 8188
rect 13443 8186 13499 8188
rect 13203 8134 13249 8186
rect 13249 8134 13259 8186
rect 13283 8134 13313 8186
rect 13313 8134 13325 8186
rect 13325 8134 13339 8186
rect 13363 8134 13377 8186
rect 13377 8134 13389 8186
rect 13389 8134 13419 8186
rect 13443 8134 13453 8186
rect 13453 8134 13499 8186
rect 13203 8132 13259 8134
rect 13283 8132 13339 8134
rect 13363 8132 13419 8134
rect 13443 8132 13499 8134
rect 10753 6554 10809 6556
rect 10833 6554 10889 6556
rect 10913 6554 10969 6556
rect 10993 6554 11049 6556
rect 10753 6502 10799 6554
rect 10799 6502 10809 6554
rect 10833 6502 10863 6554
rect 10863 6502 10875 6554
rect 10875 6502 10889 6554
rect 10913 6502 10927 6554
rect 10927 6502 10939 6554
rect 10939 6502 10969 6554
rect 10993 6502 11003 6554
rect 11003 6502 11049 6554
rect 10753 6500 10809 6502
rect 10833 6500 10889 6502
rect 10913 6500 10969 6502
rect 10993 6500 11049 6502
rect 10753 5466 10809 5468
rect 10833 5466 10889 5468
rect 10913 5466 10969 5468
rect 10993 5466 11049 5468
rect 10753 5414 10799 5466
rect 10799 5414 10809 5466
rect 10833 5414 10863 5466
rect 10863 5414 10875 5466
rect 10875 5414 10889 5466
rect 10913 5414 10927 5466
rect 10927 5414 10939 5466
rect 10939 5414 10969 5466
rect 10993 5414 11003 5466
rect 11003 5414 11049 5466
rect 10753 5412 10809 5414
rect 10833 5412 10889 5414
rect 10913 5412 10969 5414
rect 10993 5412 11049 5414
rect 10753 4378 10809 4380
rect 10833 4378 10889 4380
rect 10913 4378 10969 4380
rect 10993 4378 11049 4380
rect 10753 4326 10799 4378
rect 10799 4326 10809 4378
rect 10833 4326 10863 4378
rect 10863 4326 10875 4378
rect 10875 4326 10889 4378
rect 10913 4326 10927 4378
rect 10927 4326 10939 4378
rect 10939 4326 10969 4378
rect 10993 4326 11003 4378
rect 11003 4326 11049 4378
rect 10753 4324 10809 4326
rect 10833 4324 10889 4326
rect 10913 4324 10969 4326
rect 10993 4324 11049 4326
rect 13203 7098 13259 7100
rect 13283 7098 13339 7100
rect 13363 7098 13419 7100
rect 13443 7098 13499 7100
rect 13203 7046 13249 7098
rect 13249 7046 13259 7098
rect 13283 7046 13313 7098
rect 13313 7046 13325 7098
rect 13325 7046 13339 7098
rect 13363 7046 13377 7098
rect 13377 7046 13389 7098
rect 13389 7046 13419 7098
rect 13443 7046 13453 7098
rect 13453 7046 13499 7098
rect 13203 7044 13259 7046
rect 13283 7044 13339 7046
rect 13363 7044 13419 7046
rect 13443 7044 13499 7046
rect 15652 20698 15708 20700
rect 15732 20698 15788 20700
rect 15812 20698 15868 20700
rect 15892 20698 15948 20700
rect 15652 20646 15698 20698
rect 15698 20646 15708 20698
rect 15732 20646 15762 20698
rect 15762 20646 15774 20698
rect 15774 20646 15788 20698
rect 15812 20646 15826 20698
rect 15826 20646 15838 20698
rect 15838 20646 15868 20698
rect 15892 20646 15902 20698
rect 15902 20646 15948 20698
rect 15652 20644 15708 20646
rect 15732 20644 15788 20646
rect 15812 20644 15868 20646
rect 15892 20644 15948 20646
rect 15652 19610 15708 19612
rect 15732 19610 15788 19612
rect 15812 19610 15868 19612
rect 15892 19610 15948 19612
rect 15652 19558 15698 19610
rect 15698 19558 15708 19610
rect 15732 19558 15762 19610
rect 15762 19558 15774 19610
rect 15774 19558 15788 19610
rect 15812 19558 15826 19610
rect 15826 19558 15838 19610
rect 15838 19558 15868 19610
rect 15892 19558 15902 19610
rect 15902 19558 15948 19610
rect 15652 19556 15708 19558
rect 15732 19556 15788 19558
rect 15812 19556 15868 19558
rect 15892 19556 15948 19558
rect 15652 18522 15708 18524
rect 15732 18522 15788 18524
rect 15812 18522 15868 18524
rect 15892 18522 15948 18524
rect 15652 18470 15698 18522
rect 15698 18470 15708 18522
rect 15732 18470 15762 18522
rect 15762 18470 15774 18522
rect 15774 18470 15788 18522
rect 15812 18470 15826 18522
rect 15826 18470 15838 18522
rect 15838 18470 15868 18522
rect 15892 18470 15902 18522
rect 15902 18470 15948 18522
rect 15652 18468 15708 18470
rect 15732 18468 15788 18470
rect 15812 18468 15868 18470
rect 15892 18468 15948 18470
rect 13203 6010 13259 6012
rect 13283 6010 13339 6012
rect 13363 6010 13419 6012
rect 13443 6010 13499 6012
rect 13203 5958 13249 6010
rect 13249 5958 13259 6010
rect 13283 5958 13313 6010
rect 13313 5958 13325 6010
rect 13325 5958 13339 6010
rect 13363 5958 13377 6010
rect 13377 5958 13389 6010
rect 13389 5958 13419 6010
rect 13443 5958 13453 6010
rect 13453 5958 13499 6010
rect 13203 5956 13259 5958
rect 13283 5956 13339 5958
rect 13363 5956 13419 5958
rect 13443 5956 13499 5958
rect 13203 4922 13259 4924
rect 13283 4922 13339 4924
rect 13363 4922 13419 4924
rect 13443 4922 13499 4924
rect 13203 4870 13249 4922
rect 13249 4870 13259 4922
rect 13283 4870 13313 4922
rect 13313 4870 13325 4922
rect 13325 4870 13339 4922
rect 13363 4870 13377 4922
rect 13377 4870 13389 4922
rect 13389 4870 13419 4922
rect 13443 4870 13453 4922
rect 13453 4870 13499 4922
rect 13203 4868 13259 4870
rect 13283 4868 13339 4870
rect 13363 4868 13419 4870
rect 13443 4868 13499 4870
rect 5854 2202 5910 2204
rect 5934 2202 5990 2204
rect 6014 2202 6070 2204
rect 6094 2202 6150 2204
rect 5854 2150 5900 2202
rect 5900 2150 5910 2202
rect 5934 2150 5964 2202
rect 5964 2150 5976 2202
rect 5976 2150 5990 2202
rect 6014 2150 6028 2202
rect 6028 2150 6040 2202
rect 6040 2150 6070 2202
rect 6094 2150 6104 2202
rect 6104 2150 6150 2202
rect 5854 2148 5910 2150
rect 5934 2148 5990 2150
rect 6014 2148 6070 2150
rect 6094 2148 6150 2150
rect 10753 3290 10809 3292
rect 10833 3290 10889 3292
rect 10913 3290 10969 3292
rect 10993 3290 11049 3292
rect 10753 3238 10799 3290
rect 10799 3238 10809 3290
rect 10833 3238 10863 3290
rect 10863 3238 10875 3290
rect 10875 3238 10889 3290
rect 10913 3238 10927 3290
rect 10927 3238 10939 3290
rect 10939 3238 10969 3290
rect 10993 3238 11003 3290
rect 11003 3238 11049 3290
rect 10753 3236 10809 3238
rect 10833 3236 10889 3238
rect 10913 3236 10969 3238
rect 10993 3236 11049 3238
rect 13203 3834 13259 3836
rect 13283 3834 13339 3836
rect 13363 3834 13419 3836
rect 13443 3834 13499 3836
rect 13203 3782 13249 3834
rect 13249 3782 13259 3834
rect 13283 3782 13313 3834
rect 13313 3782 13325 3834
rect 13325 3782 13339 3834
rect 13363 3782 13377 3834
rect 13377 3782 13389 3834
rect 13389 3782 13419 3834
rect 13443 3782 13453 3834
rect 13453 3782 13499 3834
rect 13203 3780 13259 3782
rect 13283 3780 13339 3782
rect 13363 3780 13419 3782
rect 13443 3780 13499 3782
rect 13203 2746 13259 2748
rect 13283 2746 13339 2748
rect 13363 2746 13419 2748
rect 13443 2746 13499 2748
rect 13203 2694 13249 2746
rect 13249 2694 13259 2746
rect 13283 2694 13313 2746
rect 13313 2694 13325 2746
rect 13325 2694 13339 2746
rect 13363 2694 13377 2746
rect 13377 2694 13389 2746
rect 13389 2694 13419 2746
rect 13443 2694 13453 2746
rect 13453 2694 13499 2746
rect 13203 2692 13259 2694
rect 13283 2692 13339 2694
rect 13363 2692 13419 2694
rect 13443 2692 13499 2694
rect 15652 17434 15708 17436
rect 15732 17434 15788 17436
rect 15812 17434 15868 17436
rect 15892 17434 15948 17436
rect 15652 17382 15698 17434
rect 15698 17382 15708 17434
rect 15732 17382 15762 17434
rect 15762 17382 15774 17434
rect 15774 17382 15788 17434
rect 15812 17382 15826 17434
rect 15826 17382 15838 17434
rect 15838 17382 15868 17434
rect 15892 17382 15902 17434
rect 15902 17382 15948 17434
rect 15652 17380 15708 17382
rect 15732 17380 15788 17382
rect 15812 17380 15868 17382
rect 15892 17380 15948 17382
rect 18102 21242 18158 21244
rect 18182 21242 18238 21244
rect 18262 21242 18318 21244
rect 18342 21242 18398 21244
rect 18102 21190 18148 21242
rect 18148 21190 18158 21242
rect 18182 21190 18212 21242
rect 18212 21190 18224 21242
rect 18224 21190 18238 21242
rect 18262 21190 18276 21242
rect 18276 21190 18288 21242
rect 18288 21190 18318 21242
rect 18342 21190 18352 21242
rect 18352 21190 18398 21242
rect 18102 21188 18158 21190
rect 18182 21188 18238 21190
rect 18262 21188 18318 21190
rect 18342 21188 18398 21190
rect 18102 20154 18158 20156
rect 18182 20154 18238 20156
rect 18262 20154 18318 20156
rect 18342 20154 18398 20156
rect 18102 20102 18148 20154
rect 18148 20102 18158 20154
rect 18182 20102 18212 20154
rect 18212 20102 18224 20154
rect 18224 20102 18238 20154
rect 18262 20102 18276 20154
rect 18276 20102 18288 20154
rect 18288 20102 18318 20154
rect 18342 20102 18352 20154
rect 18352 20102 18398 20154
rect 18102 20100 18158 20102
rect 18182 20100 18238 20102
rect 18262 20100 18318 20102
rect 18342 20100 18398 20102
rect 18102 19066 18158 19068
rect 18182 19066 18238 19068
rect 18262 19066 18318 19068
rect 18342 19066 18398 19068
rect 18102 19014 18148 19066
rect 18148 19014 18158 19066
rect 18182 19014 18212 19066
rect 18212 19014 18224 19066
rect 18224 19014 18238 19066
rect 18262 19014 18276 19066
rect 18276 19014 18288 19066
rect 18288 19014 18318 19066
rect 18342 19014 18352 19066
rect 18352 19014 18398 19066
rect 18102 19012 18158 19014
rect 18182 19012 18238 19014
rect 18262 19012 18318 19014
rect 18342 19012 18398 19014
rect 15652 16346 15708 16348
rect 15732 16346 15788 16348
rect 15812 16346 15868 16348
rect 15892 16346 15948 16348
rect 15652 16294 15698 16346
rect 15698 16294 15708 16346
rect 15732 16294 15762 16346
rect 15762 16294 15774 16346
rect 15774 16294 15788 16346
rect 15812 16294 15826 16346
rect 15826 16294 15838 16346
rect 15838 16294 15868 16346
rect 15892 16294 15902 16346
rect 15902 16294 15948 16346
rect 15652 16292 15708 16294
rect 15732 16292 15788 16294
rect 15812 16292 15868 16294
rect 15892 16292 15948 16294
rect 18102 17978 18158 17980
rect 18182 17978 18238 17980
rect 18262 17978 18318 17980
rect 18342 17978 18398 17980
rect 18102 17926 18148 17978
rect 18148 17926 18158 17978
rect 18182 17926 18212 17978
rect 18212 17926 18224 17978
rect 18224 17926 18238 17978
rect 18262 17926 18276 17978
rect 18276 17926 18288 17978
rect 18288 17926 18318 17978
rect 18342 17926 18352 17978
rect 18352 17926 18398 17978
rect 18102 17924 18158 17926
rect 18182 17924 18238 17926
rect 18262 17924 18318 17926
rect 18342 17924 18398 17926
rect 15652 15258 15708 15260
rect 15732 15258 15788 15260
rect 15812 15258 15868 15260
rect 15892 15258 15948 15260
rect 15652 15206 15698 15258
rect 15698 15206 15708 15258
rect 15732 15206 15762 15258
rect 15762 15206 15774 15258
rect 15774 15206 15788 15258
rect 15812 15206 15826 15258
rect 15826 15206 15838 15258
rect 15838 15206 15868 15258
rect 15892 15206 15902 15258
rect 15902 15206 15948 15258
rect 15652 15204 15708 15206
rect 15732 15204 15788 15206
rect 15812 15204 15868 15206
rect 15892 15204 15948 15206
rect 15652 14170 15708 14172
rect 15732 14170 15788 14172
rect 15812 14170 15868 14172
rect 15892 14170 15948 14172
rect 15652 14118 15698 14170
rect 15698 14118 15708 14170
rect 15732 14118 15762 14170
rect 15762 14118 15774 14170
rect 15774 14118 15788 14170
rect 15812 14118 15826 14170
rect 15826 14118 15838 14170
rect 15838 14118 15868 14170
rect 15892 14118 15902 14170
rect 15902 14118 15948 14170
rect 15652 14116 15708 14118
rect 15732 14116 15788 14118
rect 15812 14116 15868 14118
rect 15892 14116 15948 14118
rect 15652 13082 15708 13084
rect 15732 13082 15788 13084
rect 15812 13082 15868 13084
rect 15892 13082 15948 13084
rect 15652 13030 15698 13082
rect 15698 13030 15708 13082
rect 15732 13030 15762 13082
rect 15762 13030 15774 13082
rect 15774 13030 15788 13082
rect 15812 13030 15826 13082
rect 15826 13030 15838 13082
rect 15838 13030 15868 13082
rect 15892 13030 15902 13082
rect 15902 13030 15948 13082
rect 15652 13028 15708 13030
rect 15732 13028 15788 13030
rect 15812 13028 15868 13030
rect 15892 13028 15948 13030
rect 15652 11994 15708 11996
rect 15732 11994 15788 11996
rect 15812 11994 15868 11996
rect 15892 11994 15948 11996
rect 15652 11942 15698 11994
rect 15698 11942 15708 11994
rect 15732 11942 15762 11994
rect 15762 11942 15774 11994
rect 15774 11942 15788 11994
rect 15812 11942 15826 11994
rect 15826 11942 15838 11994
rect 15838 11942 15868 11994
rect 15892 11942 15902 11994
rect 15902 11942 15948 11994
rect 15652 11940 15708 11942
rect 15732 11940 15788 11942
rect 15812 11940 15868 11942
rect 15892 11940 15948 11942
rect 15652 10906 15708 10908
rect 15732 10906 15788 10908
rect 15812 10906 15868 10908
rect 15892 10906 15948 10908
rect 15652 10854 15698 10906
rect 15698 10854 15708 10906
rect 15732 10854 15762 10906
rect 15762 10854 15774 10906
rect 15774 10854 15788 10906
rect 15812 10854 15826 10906
rect 15826 10854 15838 10906
rect 15838 10854 15868 10906
rect 15892 10854 15902 10906
rect 15902 10854 15948 10906
rect 15652 10852 15708 10854
rect 15732 10852 15788 10854
rect 15812 10852 15868 10854
rect 15892 10852 15948 10854
rect 15652 9818 15708 9820
rect 15732 9818 15788 9820
rect 15812 9818 15868 9820
rect 15892 9818 15948 9820
rect 15652 9766 15698 9818
rect 15698 9766 15708 9818
rect 15732 9766 15762 9818
rect 15762 9766 15774 9818
rect 15774 9766 15788 9818
rect 15812 9766 15826 9818
rect 15826 9766 15838 9818
rect 15838 9766 15868 9818
rect 15892 9766 15902 9818
rect 15902 9766 15948 9818
rect 15652 9764 15708 9766
rect 15732 9764 15788 9766
rect 15812 9764 15868 9766
rect 15892 9764 15948 9766
rect 15652 8730 15708 8732
rect 15732 8730 15788 8732
rect 15812 8730 15868 8732
rect 15892 8730 15948 8732
rect 15652 8678 15698 8730
rect 15698 8678 15708 8730
rect 15732 8678 15762 8730
rect 15762 8678 15774 8730
rect 15774 8678 15788 8730
rect 15812 8678 15826 8730
rect 15826 8678 15838 8730
rect 15838 8678 15868 8730
rect 15892 8678 15902 8730
rect 15902 8678 15948 8730
rect 15652 8676 15708 8678
rect 15732 8676 15788 8678
rect 15812 8676 15868 8678
rect 15892 8676 15948 8678
rect 15652 7642 15708 7644
rect 15732 7642 15788 7644
rect 15812 7642 15868 7644
rect 15892 7642 15948 7644
rect 15652 7590 15698 7642
rect 15698 7590 15708 7642
rect 15732 7590 15762 7642
rect 15762 7590 15774 7642
rect 15774 7590 15788 7642
rect 15812 7590 15826 7642
rect 15826 7590 15838 7642
rect 15838 7590 15868 7642
rect 15892 7590 15902 7642
rect 15902 7590 15948 7642
rect 15652 7588 15708 7590
rect 15732 7588 15788 7590
rect 15812 7588 15868 7590
rect 15892 7588 15948 7590
rect 15652 6554 15708 6556
rect 15732 6554 15788 6556
rect 15812 6554 15868 6556
rect 15892 6554 15948 6556
rect 15652 6502 15698 6554
rect 15698 6502 15708 6554
rect 15732 6502 15762 6554
rect 15762 6502 15774 6554
rect 15774 6502 15788 6554
rect 15812 6502 15826 6554
rect 15826 6502 15838 6554
rect 15838 6502 15868 6554
rect 15892 6502 15902 6554
rect 15902 6502 15948 6554
rect 15652 6500 15708 6502
rect 15732 6500 15788 6502
rect 15812 6500 15868 6502
rect 15892 6500 15948 6502
rect 15652 5466 15708 5468
rect 15732 5466 15788 5468
rect 15812 5466 15868 5468
rect 15892 5466 15948 5468
rect 15652 5414 15698 5466
rect 15698 5414 15708 5466
rect 15732 5414 15762 5466
rect 15762 5414 15774 5466
rect 15774 5414 15788 5466
rect 15812 5414 15826 5466
rect 15826 5414 15838 5466
rect 15838 5414 15868 5466
rect 15892 5414 15902 5466
rect 15902 5414 15948 5466
rect 15652 5412 15708 5414
rect 15732 5412 15788 5414
rect 15812 5412 15868 5414
rect 15892 5412 15948 5414
rect 15652 4378 15708 4380
rect 15732 4378 15788 4380
rect 15812 4378 15868 4380
rect 15892 4378 15948 4380
rect 15652 4326 15698 4378
rect 15698 4326 15708 4378
rect 15732 4326 15762 4378
rect 15762 4326 15774 4378
rect 15774 4326 15788 4378
rect 15812 4326 15826 4378
rect 15826 4326 15838 4378
rect 15838 4326 15868 4378
rect 15892 4326 15902 4378
rect 15902 4326 15948 4378
rect 15652 4324 15708 4326
rect 15732 4324 15788 4326
rect 15812 4324 15868 4326
rect 15892 4324 15948 4326
rect 15652 3290 15708 3292
rect 15732 3290 15788 3292
rect 15812 3290 15868 3292
rect 15892 3290 15948 3292
rect 15652 3238 15698 3290
rect 15698 3238 15708 3290
rect 15732 3238 15762 3290
rect 15762 3238 15774 3290
rect 15774 3238 15788 3290
rect 15812 3238 15826 3290
rect 15826 3238 15838 3290
rect 15838 3238 15868 3290
rect 15892 3238 15902 3290
rect 15902 3238 15948 3290
rect 15652 3236 15708 3238
rect 15732 3236 15788 3238
rect 15812 3236 15868 3238
rect 15892 3236 15948 3238
rect 18102 16890 18158 16892
rect 18182 16890 18238 16892
rect 18262 16890 18318 16892
rect 18342 16890 18398 16892
rect 18102 16838 18148 16890
rect 18148 16838 18158 16890
rect 18182 16838 18212 16890
rect 18212 16838 18224 16890
rect 18224 16838 18238 16890
rect 18262 16838 18276 16890
rect 18276 16838 18288 16890
rect 18288 16838 18318 16890
rect 18342 16838 18352 16890
rect 18352 16838 18398 16890
rect 18102 16836 18158 16838
rect 18182 16836 18238 16838
rect 18262 16836 18318 16838
rect 18342 16836 18398 16838
rect 18102 15802 18158 15804
rect 18182 15802 18238 15804
rect 18262 15802 18318 15804
rect 18342 15802 18398 15804
rect 18102 15750 18148 15802
rect 18148 15750 18158 15802
rect 18182 15750 18212 15802
rect 18212 15750 18224 15802
rect 18224 15750 18238 15802
rect 18262 15750 18276 15802
rect 18276 15750 18288 15802
rect 18288 15750 18318 15802
rect 18342 15750 18352 15802
rect 18352 15750 18398 15802
rect 18102 15748 18158 15750
rect 18182 15748 18238 15750
rect 18262 15748 18318 15750
rect 18342 15748 18398 15750
rect 18102 14714 18158 14716
rect 18182 14714 18238 14716
rect 18262 14714 18318 14716
rect 18342 14714 18398 14716
rect 18102 14662 18148 14714
rect 18148 14662 18158 14714
rect 18182 14662 18212 14714
rect 18212 14662 18224 14714
rect 18224 14662 18238 14714
rect 18262 14662 18276 14714
rect 18276 14662 18288 14714
rect 18288 14662 18318 14714
rect 18342 14662 18352 14714
rect 18352 14662 18398 14714
rect 18102 14660 18158 14662
rect 18182 14660 18238 14662
rect 18262 14660 18318 14662
rect 18342 14660 18398 14662
rect 18102 13626 18158 13628
rect 18182 13626 18238 13628
rect 18262 13626 18318 13628
rect 18342 13626 18398 13628
rect 18102 13574 18148 13626
rect 18148 13574 18158 13626
rect 18182 13574 18212 13626
rect 18212 13574 18224 13626
rect 18224 13574 18238 13626
rect 18262 13574 18276 13626
rect 18276 13574 18288 13626
rect 18288 13574 18318 13626
rect 18342 13574 18352 13626
rect 18352 13574 18398 13626
rect 18102 13572 18158 13574
rect 18182 13572 18238 13574
rect 18262 13572 18318 13574
rect 18342 13572 18398 13574
rect 18102 12538 18158 12540
rect 18182 12538 18238 12540
rect 18262 12538 18318 12540
rect 18342 12538 18398 12540
rect 18102 12486 18148 12538
rect 18148 12486 18158 12538
rect 18182 12486 18212 12538
rect 18212 12486 18224 12538
rect 18224 12486 18238 12538
rect 18262 12486 18276 12538
rect 18276 12486 18288 12538
rect 18288 12486 18318 12538
rect 18342 12486 18352 12538
rect 18352 12486 18398 12538
rect 18102 12484 18158 12486
rect 18182 12484 18238 12486
rect 18262 12484 18318 12486
rect 18342 12484 18398 12486
rect 18102 11450 18158 11452
rect 18182 11450 18238 11452
rect 18262 11450 18318 11452
rect 18342 11450 18398 11452
rect 18102 11398 18148 11450
rect 18148 11398 18158 11450
rect 18182 11398 18212 11450
rect 18212 11398 18224 11450
rect 18224 11398 18238 11450
rect 18262 11398 18276 11450
rect 18276 11398 18288 11450
rect 18288 11398 18318 11450
rect 18342 11398 18352 11450
rect 18352 11398 18398 11450
rect 18102 11396 18158 11398
rect 18182 11396 18238 11398
rect 18262 11396 18318 11398
rect 18342 11396 18398 11398
rect 19246 15000 19302 15056
rect 18102 10362 18158 10364
rect 18182 10362 18238 10364
rect 18262 10362 18318 10364
rect 18342 10362 18398 10364
rect 18102 10310 18148 10362
rect 18148 10310 18158 10362
rect 18182 10310 18212 10362
rect 18212 10310 18224 10362
rect 18224 10310 18238 10362
rect 18262 10310 18276 10362
rect 18276 10310 18288 10362
rect 18288 10310 18318 10362
rect 18342 10310 18352 10362
rect 18352 10310 18398 10362
rect 18102 10308 18158 10310
rect 18182 10308 18238 10310
rect 18262 10308 18318 10310
rect 18342 10308 18398 10310
rect 18102 9274 18158 9276
rect 18182 9274 18238 9276
rect 18262 9274 18318 9276
rect 18342 9274 18398 9276
rect 18102 9222 18148 9274
rect 18148 9222 18158 9274
rect 18182 9222 18212 9274
rect 18212 9222 18224 9274
rect 18224 9222 18238 9274
rect 18262 9222 18276 9274
rect 18276 9222 18288 9274
rect 18288 9222 18318 9274
rect 18342 9222 18352 9274
rect 18352 9222 18398 9274
rect 18102 9220 18158 9222
rect 18182 9220 18238 9222
rect 18262 9220 18318 9222
rect 18342 9220 18398 9222
rect 18102 8186 18158 8188
rect 18182 8186 18238 8188
rect 18262 8186 18318 8188
rect 18342 8186 18398 8188
rect 18102 8134 18148 8186
rect 18148 8134 18158 8186
rect 18182 8134 18212 8186
rect 18212 8134 18224 8186
rect 18224 8134 18238 8186
rect 18262 8134 18276 8186
rect 18276 8134 18288 8186
rect 18288 8134 18318 8186
rect 18342 8134 18352 8186
rect 18352 8134 18398 8186
rect 18102 8132 18158 8134
rect 18182 8132 18238 8134
rect 18262 8132 18318 8134
rect 18342 8132 18398 8134
rect 18102 7098 18158 7100
rect 18182 7098 18238 7100
rect 18262 7098 18318 7100
rect 18342 7098 18398 7100
rect 18102 7046 18148 7098
rect 18148 7046 18158 7098
rect 18182 7046 18212 7098
rect 18212 7046 18224 7098
rect 18224 7046 18238 7098
rect 18262 7046 18276 7098
rect 18276 7046 18288 7098
rect 18288 7046 18318 7098
rect 18342 7046 18352 7098
rect 18352 7046 18398 7098
rect 18102 7044 18158 7046
rect 18182 7044 18238 7046
rect 18262 7044 18318 7046
rect 18342 7044 18398 7046
rect 18102 6010 18158 6012
rect 18182 6010 18238 6012
rect 18262 6010 18318 6012
rect 18342 6010 18398 6012
rect 18102 5958 18148 6010
rect 18148 5958 18158 6010
rect 18182 5958 18212 6010
rect 18212 5958 18224 6010
rect 18224 5958 18238 6010
rect 18262 5958 18276 6010
rect 18276 5958 18288 6010
rect 18288 5958 18318 6010
rect 18342 5958 18352 6010
rect 18352 5958 18398 6010
rect 18102 5956 18158 5958
rect 18182 5956 18238 5958
rect 18262 5956 18318 5958
rect 18342 5956 18398 5958
rect 18102 4922 18158 4924
rect 18182 4922 18238 4924
rect 18262 4922 18318 4924
rect 18342 4922 18398 4924
rect 18102 4870 18148 4922
rect 18148 4870 18158 4922
rect 18182 4870 18212 4922
rect 18212 4870 18224 4922
rect 18224 4870 18238 4922
rect 18262 4870 18276 4922
rect 18276 4870 18288 4922
rect 18288 4870 18318 4922
rect 18342 4870 18352 4922
rect 18352 4870 18398 4922
rect 18102 4868 18158 4870
rect 18182 4868 18238 4870
rect 18262 4868 18318 4870
rect 18342 4868 18398 4870
rect 18102 3834 18158 3836
rect 18182 3834 18238 3836
rect 18262 3834 18318 3836
rect 18342 3834 18398 3836
rect 18102 3782 18148 3834
rect 18148 3782 18158 3834
rect 18182 3782 18212 3834
rect 18212 3782 18224 3834
rect 18224 3782 18238 3834
rect 18262 3782 18276 3834
rect 18276 3782 18288 3834
rect 18288 3782 18318 3834
rect 18342 3782 18352 3834
rect 18352 3782 18398 3834
rect 18102 3780 18158 3782
rect 18182 3780 18238 3782
rect 18262 3780 18318 3782
rect 18342 3780 18398 3782
rect 18102 2746 18158 2748
rect 18182 2746 18238 2748
rect 18262 2746 18318 2748
rect 18342 2746 18398 2748
rect 18102 2694 18148 2746
rect 18148 2694 18158 2746
rect 18182 2694 18212 2746
rect 18212 2694 18224 2746
rect 18224 2694 18238 2746
rect 18262 2694 18276 2746
rect 18276 2694 18288 2746
rect 18288 2694 18318 2746
rect 18342 2694 18352 2746
rect 18352 2694 18398 2746
rect 18102 2692 18158 2694
rect 18182 2692 18238 2694
rect 18262 2692 18318 2694
rect 18342 2692 18398 2694
rect 20551 20698 20607 20700
rect 20631 20698 20687 20700
rect 20711 20698 20767 20700
rect 20791 20698 20847 20700
rect 20551 20646 20597 20698
rect 20597 20646 20607 20698
rect 20631 20646 20661 20698
rect 20661 20646 20673 20698
rect 20673 20646 20687 20698
rect 20711 20646 20725 20698
rect 20725 20646 20737 20698
rect 20737 20646 20767 20698
rect 20791 20646 20801 20698
rect 20801 20646 20847 20698
rect 20551 20644 20607 20646
rect 20631 20644 20687 20646
rect 20711 20644 20767 20646
rect 20791 20644 20847 20646
rect 20350 19896 20406 19952
rect 20551 19610 20607 19612
rect 20631 19610 20687 19612
rect 20711 19610 20767 19612
rect 20791 19610 20847 19612
rect 20551 19558 20597 19610
rect 20597 19558 20607 19610
rect 20631 19558 20661 19610
rect 20661 19558 20673 19610
rect 20673 19558 20687 19610
rect 20711 19558 20725 19610
rect 20725 19558 20737 19610
rect 20737 19558 20767 19610
rect 20791 19558 20801 19610
rect 20801 19558 20847 19610
rect 20551 19556 20607 19558
rect 20631 19556 20687 19558
rect 20711 19556 20767 19558
rect 20791 19556 20847 19558
rect 20551 18522 20607 18524
rect 20631 18522 20687 18524
rect 20711 18522 20767 18524
rect 20791 18522 20847 18524
rect 20551 18470 20597 18522
rect 20597 18470 20607 18522
rect 20631 18470 20661 18522
rect 20661 18470 20673 18522
rect 20673 18470 20687 18522
rect 20711 18470 20725 18522
rect 20725 18470 20737 18522
rect 20737 18470 20767 18522
rect 20791 18470 20801 18522
rect 20801 18470 20847 18522
rect 20551 18468 20607 18470
rect 20631 18468 20687 18470
rect 20711 18468 20767 18470
rect 20791 18468 20847 18470
rect 20258 18264 20314 18320
rect 20551 17434 20607 17436
rect 20631 17434 20687 17436
rect 20711 17434 20767 17436
rect 20791 17434 20847 17436
rect 20551 17382 20597 17434
rect 20597 17382 20607 17434
rect 20631 17382 20661 17434
rect 20661 17382 20673 17434
rect 20673 17382 20687 17434
rect 20711 17382 20725 17434
rect 20725 17382 20737 17434
rect 20737 17382 20767 17434
rect 20791 17382 20801 17434
rect 20801 17382 20847 17434
rect 20551 17380 20607 17382
rect 20631 17380 20687 17382
rect 20711 17380 20767 17382
rect 20791 17380 20847 17382
rect 20258 16632 20314 16688
rect 20166 13404 20168 13424
rect 20168 13404 20220 13424
rect 20220 13404 20222 13424
rect 20166 13368 20222 13404
rect 20166 11736 20222 11792
rect 20166 10140 20168 10160
rect 20168 10140 20220 10160
rect 20220 10140 20222 10160
rect 20166 10104 20222 10140
rect 20166 8472 20222 8528
rect 20166 6840 20222 6896
rect 20258 5208 20314 5264
rect 20258 3612 20260 3632
rect 20260 3612 20312 3632
rect 20312 3612 20314 3632
rect 20258 3576 20314 3612
rect 10753 2202 10809 2204
rect 10833 2202 10889 2204
rect 10913 2202 10969 2204
rect 10993 2202 11049 2204
rect 10753 2150 10799 2202
rect 10799 2150 10809 2202
rect 10833 2150 10863 2202
rect 10863 2150 10875 2202
rect 10875 2150 10889 2202
rect 10913 2150 10927 2202
rect 10927 2150 10939 2202
rect 10939 2150 10969 2202
rect 10993 2150 11003 2202
rect 11003 2150 11049 2202
rect 10753 2148 10809 2150
rect 10833 2148 10889 2150
rect 10913 2148 10969 2150
rect 10993 2148 11049 2150
rect 15652 2202 15708 2204
rect 15732 2202 15788 2204
rect 15812 2202 15868 2204
rect 15892 2202 15948 2204
rect 15652 2150 15698 2202
rect 15698 2150 15708 2202
rect 15732 2150 15762 2202
rect 15762 2150 15774 2202
rect 15774 2150 15788 2202
rect 15812 2150 15826 2202
rect 15826 2150 15838 2202
rect 15838 2150 15868 2202
rect 15892 2150 15902 2202
rect 15902 2150 15948 2202
rect 15652 2148 15708 2150
rect 15732 2148 15788 2150
rect 15812 2148 15868 2150
rect 15892 2148 15948 2150
rect 20551 16346 20607 16348
rect 20631 16346 20687 16348
rect 20711 16346 20767 16348
rect 20791 16346 20847 16348
rect 20551 16294 20597 16346
rect 20597 16294 20607 16346
rect 20631 16294 20661 16346
rect 20661 16294 20673 16346
rect 20673 16294 20687 16346
rect 20711 16294 20725 16346
rect 20725 16294 20737 16346
rect 20737 16294 20767 16346
rect 20791 16294 20801 16346
rect 20801 16294 20847 16346
rect 20551 16292 20607 16294
rect 20631 16292 20687 16294
rect 20711 16292 20767 16294
rect 20791 16292 20847 16294
rect 20551 15258 20607 15260
rect 20631 15258 20687 15260
rect 20711 15258 20767 15260
rect 20791 15258 20847 15260
rect 20551 15206 20597 15258
rect 20597 15206 20607 15258
rect 20631 15206 20661 15258
rect 20661 15206 20673 15258
rect 20673 15206 20687 15258
rect 20711 15206 20725 15258
rect 20725 15206 20737 15258
rect 20737 15206 20767 15258
rect 20791 15206 20801 15258
rect 20801 15206 20847 15258
rect 20551 15204 20607 15206
rect 20631 15204 20687 15206
rect 20711 15204 20767 15206
rect 20791 15204 20847 15206
rect 20551 14170 20607 14172
rect 20631 14170 20687 14172
rect 20711 14170 20767 14172
rect 20791 14170 20847 14172
rect 20551 14118 20597 14170
rect 20597 14118 20607 14170
rect 20631 14118 20661 14170
rect 20661 14118 20673 14170
rect 20673 14118 20687 14170
rect 20711 14118 20725 14170
rect 20725 14118 20737 14170
rect 20737 14118 20767 14170
rect 20791 14118 20801 14170
rect 20801 14118 20847 14170
rect 20551 14116 20607 14118
rect 20631 14116 20687 14118
rect 20711 14116 20767 14118
rect 20791 14116 20847 14118
rect 20551 13082 20607 13084
rect 20631 13082 20687 13084
rect 20711 13082 20767 13084
rect 20791 13082 20847 13084
rect 20551 13030 20597 13082
rect 20597 13030 20607 13082
rect 20631 13030 20661 13082
rect 20661 13030 20673 13082
rect 20673 13030 20687 13082
rect 20711 13030 20725 13082
rect 20725 13030 20737 13082
rect 20737 13030 20767 13082
rect 20791 13030 20801 13082
rect 20801 13030 20847 13082
rect 20551 13028 20607 13030
rect 20631 13028 20687 13030
rect 20711 13028 20767 13030
rect 20791 13028 20847 13030
rect 20551 11994 20607 11996
rect 20631 11994 20687 11996
rect 20711 11994 20767 11996
rect 20791 11994 20847 11996
rect 20551 11942 20597 11994
rect 20597 11942 20607 11994
rect 20631 11942 20661 11994
rect 20661 11942 20673 11994
rect 20673 11942 20687 11994
rect 20711 11942 20725 11994
rect 20725 11942 20737 11994
rect 20737 11942 20767 11994
rect 20791 11942 20801 11994
rect 20801 11942 20847 11994
rect 20551 11940 20607 11942
rect 20631 11940 20687 11942
rect 20711 11940 20767 11942
rect 20791 11940 20847 11942
rect 20551 10906 20607 10908
rect 20631 10906 20687 10908
rect 20711 10906 20767 10908
rect 20791 10906 20847 10908
rect 20551 10854 20597 10906
rect 20597 10854 20607 10906
rect 20631 10854 20661 10906
rect 20661 10854 20673 10906
rect 20673 10854 20687 10906
rect 20711 10854 20725 10906
rect 20725 10854 20737 10906
rect 20737 10854 20767 10906
rect 20791 10854 20801 10906
rect 20801 10854 20847 10906
rect 20551 10852 20607 10854
rect 20631 10852 20687 10854
rect 20711 10852 20767 10854
rect 20791 10852 20847 10854
rect 20551 9818 20607 9820
rect 20631 9818 20687 9820
rect 20711 9818 20767 9820
rect 20791 9818 20847 9820
rect 20551 9766 20597 9818
rect 20597 9766 20607 9818
rect 20631 9766 20661 9818
rect 20661 9766 20673 9818
rect 20673 9766 20687 9818
rect 20711 9766 20725 9818
rect 20725 9766 20737 9818
rect 20737 9766 20767 9818
rect 20791 9766 20801 9818
rect 20801 9766 20847 9818
rect 20551 9764 20607 9766
rect 20631 9764 20687 9766
rect 20711 9764 20767 9766
rect 20791 9764 20847 9766
rect 20551 8730 20607 8732
rect 20631 8730 20687 8732
rect 20711 8730 20767 8732
rect 20791 8730 20847 8732
rect 20551 8678 20597 8730
rect 20597 8678 20607 8730
rect 20631 8678 20661 8730
rect 20661 8678 20673 8730
rect 20673 8678 20687 8730
rect 20711 8678 20725 8730
rect 20725 8678 20737 8730
rect 20737 8678 20767 8730
rect 20791 8678 20801 8730
rect 20801 8678 20847 8730
rect 20551 8676 20607 8678
rect 20631 8676 20687 8678
rect 20711 8676 20767 8678
rect 20791 8676 20847 8678
rect 20551 7642 20607 7644
rect 20631 7642 20687 7644
rect 20711 7642 20767 7644
rect 20791 7642 20847 7644
rect 20551 7590 20597 7642
rect 20597 7590 20607 7642
rect 20631 7590 20661 7642
rect 20661 7590 20673 7642
rect 20673 7590 20687 7642
rect 20711 7590 20725 7642
rect 20725 7590 20737 7642
rect 20737 7590 20767 7642
rect 20791 7590 20801 7642
rect 20801 7590 20847 7642
rect 20551 7588 20607 7590
rect 20631 7588 20687 7590
rect 20711 7588 20767 7590
rect 20791 7588 20847 7590
rect 20551 6554 20607 6556
rect 20631 6554 20687 6556
rect 20711 6554 20767 6556
rect 20791 6554 20847 6556
rect 20551 6502 20597 6554
rect 20597 6502 20607 6554
rect 20631 6502 20661 6554
rect 20661 6502 20673 6554
rect 20673 6502 20687 6554
rect 20711 6502 20725 6554
rect 20725 6502 20737 6554
rect 20737 6502 20767 6554
rect 20791 6502 20801 6554
rect 20801 6502 20847 6554
rect 20551 6500 20607 6502
rect 20631 6500 20687 6502
rect 20711 6500 20767 6502
rect 20791 6500 20847 6502
rect 20551 5466 20607 5468
rect 20631 5466 20687 5468
rect 20711 5466 20767 5468
rect 20791 5466 20847 5468
rect 20551 5414 20597 5466
rect 20597 5414 20607 5466
rect 20631 5414 20661 5466
rect 20661 5414 20673 5466
rect 20673 5414 20687 5466
rect 20711 5414 20725 5466
rect 20725 5414 20737 5466
rect 20737 5414 20767 5466
rect 20791 5414 20801 5466
rect 20801 5414 20847 5466
rect 20551 5412 20607 5414
rect 20631 5412 20687 5414
rect 20711 5412 20767 5414
rect 20791 5412 20847 5414
rect 20551 4378 20607 4380
rect 20631 4378 20687 4380
rect 20711 4378 20767 4380
rect 20791 4378 20847 4380
rect 20551 4326 20597 4378
rect 20597 4326 20607 4378
rect 20631 4326 20661 4378
rect 20661 4326 20673 4378
rect 20673 4326 20687 4378
rect 20711 4326 20725 4378
rect 20725 4326 20737 4378
rect 20737 4326 20767 4378
rect 20791 4326 20801 4378
rect 20801 4326 20847 4378
rect 20551 4324 20607 4326
rect 20631 4324 20687 4326
rect 20711 4324 20767 4326
rect 20791 4324 20847 4326
rect 20551 3290 20607 3292
rect 20631 3290 20687 3292
rect 20711 3290 20767 3292
rect 20791 3290 20847 3292
rect 20551 3238 20597 3290
rect 20597 3238 20607 3290
rect 20631 3238 20661 3290
rect 20661 3238 20673 3290
rect 20673 3238 20687 3290
rect 20711 3238 20725 3290
rect 20725 3238 20737 3290
rect 20737 3238 20767 3290
rect 20791 3238 20801 3290
rect 20801 3238 20847 3290
rect 20551 3236 20607 3238
rect 20631 3236 20687 3238
rect 20711 3236 20767 3238
rect 20791 3236 20847 3238
rect 20551 2202 20607 2204
rect 20631 2202 20687 2204
rect 20711 2202 20767 2204
rect 20791 2202 20847 2204
rect 20551 2150 20597 2202
rect 20597 2150 20607 2202
rect 20631 2150 20661 2202
rect 20661 2150 20673 2202
rect 20673 2150 20687 2202
rect 20711 2150 20725 2202
rect 20725 2150 20737 2202
rect 20737 2150 20767 2202
rect 20791 2150 20801 2202
rect 20801 2150 20847 2202
rect 20551 2148 20607 2150
rect 20631 2148 20687 2150
rect 20711 2148 20767 2150
rect 20791 2148 20847 2150
rect 20166 1944 20222 2000
<< metal3 >>
rect 5844 21792 6160 21793
rect 5844 21728 5850 21792
rect 5914 21728 5930 21792
rect 5994 21728 6010 21792
rect 6074 21728 6090 21792
rect 6154 21728 6160 21792
rect 5844 21727 6160 21728
rect 10743 21792 11059 21793
rect 10743 21728 10749 21792
rect 10813 21728 10829 21792
rect 10893 21728 10909 21792
rect 10973 21728 10989 21792
rect 11053 21728 11059 21792
rect 10743 21727 11059 21728
rect 15642 21792 15958 21793
rect 15642 21728 15648 21792
rect 15712 21728 15728 21792
rect 15792 21728 15808 21792
rect 15872 21728 15888 21792
rect 15952 21728 15958 21792
rect 15642 21727 15958 21728
rect 20541 21792 20857 21793
rect 20541 21728 20547 21792
rect 20611 21728 20627 21792
rect 20691 21728 20707 21792
rect 20771 21728 20787 21792
rect 20851 21728 20857 21792
rect 20541 21727 20857 21728
rect 19609 21586 19675 21589
rect 21080 21586 21880 21616
rect 19609 21584 21880 21586
rect 19609 21528 19614 21584
rect 19670 21528 21880 21584
rect 19609 21526 21880 21528
rect 19609 21523 19675 21526
rect 21080 21496 21880 21526
rect 0 21314 800 21344
rect 1301 21314 1367 21317
rect 0 21312 1367 21314
rect 0 21256 1306 21312
rect 1362 21256 1367 21312
rect 0 21254 1367 21256
rect 0 21224 800 21254
rect 1301 21251 1367 21254
rect 3395 21248 3711 21249
rect 3395 21184 3401 21248
rect 3465 21184 3481 21248
rect 3545 21184 3561 21248
rect 3625 21184 3641 21248
rect 3705 21184 3711 21248
rect 3395 21183 3711 21184
rect 8294 21248 8610 21249
rect 8294 21184 8300 21248
rect 8364 21184 8380 21248
rect 8444 21184 8460 21248
rect 8524 21184 8540 21248
rect 8604 21184 8610 21248
rect 8294 21183 8610 21184
rect 13193 21248 13509 21249
rect 13193 21184 13199 21248
rect 13263 21184 13279 21248
rect 13343 21184 13359 21248
rect 13423 21184 13439 21248
rect 13503 21184 13509 21248
rect 13193 21183 13509 21184
rect 18092 21248 18408 21249
rect 18092 21184 18098 21248
rect 18162 21184 18178 21248
rect 18242 21184 18258 21248
rect 18322 21184 18338 21248
rect 18402 21184 18408 21248
rect 18092 21183 18408 21184
rect 5844 20704 6160 20705
rect 5844 20640 5850 20704
rect 5914 20640 5930 20704
rect 5994 20640 6010 20704
rect 6074 20640 6090 20704
rect 6154 20640 6160 20704
rect 5844 20639 6160 20640
rect 10743 20704 11059 20705
rect 10743 20640 10749 20704
rect 10813 20640 10829 20704
rect 10893 20640 10909 20704
rect 10973 20640 10989 20704
rect 11053 20640 11059 20704
rect 10743 20639 11059 20640
rect 15642 20704 15958 20705
rect 15642 20640 15648 20704
rect 15712 20640 15728 20704
rect 15792 20640 15808 20704
rect 15872 20640 15888 20704
rect 15952 20640 15958 20704
rect 15642 20639 15958 20640
rect 20541 20704 20857 20705
rect 20541 20640 20547 20704
rect 20611 20640 20627 20704
rect 20691 20640 20707 20704
rect 20771 20640 20787 20704
rect 20851 20640 20857 20704
rect 20541 20639 20857 20640
rect 3395 20160 3711 20161
rect 3395 20096 3401 20160
rect 3465 20096 3481 20160
rect 3545 20096 3561 20160
rect 3625 20096 3641 20160
rect 3705 20096 3711 20160
rect 3395 20095 3711 20096
rect 8294 20160 8610 20161
rect 8294 20096 8300 20160
rect 8364 20096 8380 20160
rect 8444 20096 8460 20160
rect 8524 20096 8540 20160
rect 8604 20096 8610 20160
rect 8294 20095 8610 20096
rect 13193 20160 13509 20161
rect 13193 20096 13199 20160
rect 13263 20096 13279 20160
rect 13343 20096 13359 20160
rect 13423 20096 13439 20160
rect 13503 20096 13509 20160
rect 13193 20095 13509 20096
rect 18092 20160 18408 20161
rect 18092 20096 18098 20160
rect 18162 20096 18178 20160
rect 18242 20096 18258 20160
rect 18322 20096 18338 20160
rect 18402 20096 18408 20160
rect 18092 20095 18408 20096
rect 20345 19954 20411 19957
rect 21080 19954 21880 19984
rect 20345 19952 21880 19954
rect 20345 19896 20350 19952
rect 20406 19896 21880 19952
rect 20345 19894 21880 19896
rect 20345 19891 20411 19894
rect 21080 19864 21880 19894
rect 5844 19616 6160 19617
rect 5844 19552 5850 19616
rect 5914 19552 5930 19616
rect 5994 19552 6010 19616
rect 6074 19552 6090 19616
rect 6154 19552 6160 19616
rect 5844 19551 6160 19552
rect 10743 19616 11059 19617
rect 10743 19552 10749 19616
rect 10813 19552 10829 19616
rect 10893 19552 10909 19616
rect 10973 19552 10989 19616
rect 11053 19552 11059 19616
rect 10743 19551 11059 19552
rect 15642 19616 15958 19617
rect 15642 19552 15648 19616
rect 15712 19552 15728 19616
rect 15792 19552 15808 19616
rect 15872 19552 15888 19616
rect 15952 19552 15958 19616
rect 15642 19551 15958 19552
rect 20541 19616 20857 19617
rect 20541 19552 20547 19616
rect 20611 19552 20627 19616
rect 20691 19552 20707 19616
rect 20771 19552 20787 19616
rect 20851 19552 20857 19616
rect 20541 19551 20857 19552
rect 3395 19072 3711 19073
rect 3395 19008 3401 19072
rect 3465 19008 3481 19072
rect 3545 19008 3561 19072
rect 3625 19008 3641 19072
rect 3705 19008 3711 19072
rect 3395 19007 3711 19008
rect 8294 19072 8610 19073
rect 8294 19008 8300 19072
rect 8364 19008 8380 19072
rect 8444 19008 8460 19072
rect 8524 19008 8540 19072
rect 8604 19008 8610 19072
rect 8294 19007 8610 19008
rect 13193 19072 13509 19073
rect 13193 19008 13199 19072
rect 13263 19008 13279 19072
rect 13343 19008 13359 19072
rect 13423 19008 13439 19072
rect 13503 19008 13509 19072
rect 13193 19007 13509 19008
rect 18092 19072 18408 19073
rect 18092 19008 18098 19072
rect 18162 19008 18178 19072
rect 18242 19008 18258 19072
rect 18322 19008 18338 19072
rect 18402 19008 18408 19072
rect 18092 19007 18408 19008
rect 5844 18528 6160 18529
rect 5844 18464 5850 18528
rect 5914 18464 5930 18528
rect 5994 18464 6010 18528
rect 6074 18464 6090 18528
rect 6154 18464 6160 18528
rect 5844 18463 6160 18464
rect 10743 18528 11059 18529
rect 10743 18464 10749 18528
rect 10813 18464 10829 18528
rect 10893 18464 10909 18528
rect 10973 18464 10989 18528
rect 11053 18464 11059 18528
rect 10743 18463 11059 18464
rect 15642 18528 15958 18529
rect 15642 18464 15648 18528
rect 15712 18464 15728 18528
rect 15792 18464 15808 18528
rect 15872 18464 15888 18528
rect 15952 18464 15958 18528
rect 15642 18463 15958 18464
rect 20541 18528 20857 18529
rect 20541 18464 20547 18528
rect 20611 18464 20627 18528
rect 20691 18464 20707 18528
rect 20771 18464 20787 18528
rect 20851 18464 20857 18528
rect 20541 18463 20857 18464
rect 20253 18322 20319 18325
rect 21080 18322 21880 18352
rect 20253 18320 21880 18322
rect 20253 18264 20258 18320
rect 20314 18264 21880 18320
rect 20253 18262 21880 18264
rect 20253 18259 20319 18262
rect 21080 18232 21880 18262
rect 3395 17984 3711 17985
rect 3395 17920 3401 17984
rect 3465 17920 3481 17984
rect 3545 17920 3561 17984
rect 3625 17920 3641 17984
rect 3705 17920 3711 17984
rect 3395 17919 3711 17920
rect 8294 17984 8610 17985
rect 8294 17920 8300 17984
rect 8364 17920 8380 17984
rect 8444 17920 8460 17984
rect 8524 17920 8540 17984
rect 8604 17920 8610 17984
rect 8294 17919 8610 17920
rect 13193 17984 13509 17985
rect 13193 17920 13199 17984
rect 13263 17920 13279 17984
rect 13343 17920 13359 17984
rect 13423 17920 13439 17984
rect 13503 17920 13509 17984
rect 13193 17919 13509 17920
rect 18092 17984 18408 17985
rect 18092 17920 18098 17984
rect 18162 17920 18178 17984
rect 18242 17920 18258 17984
rect 18322 17920 18338 17984
rect 18402 17920 18408 17984
rect 18092 17919 18408 17920
rect 0 17416 800 17536
rect 5844 17440 6160 17441
rect 5844 17376 5850 17440
rect 5914 17376 5930 17440
rect 5994 17376 6010 17440
rect 6074 17376 6090 17440
rect 6154 17376 6160 17440
rect 5844 17375 6160 17376
rect 10743 17440 11059 17441
rect 10743 17376 10749 17440
rect 10813 17376 10829 17440
rect 10893 17376 10909 17440
rect 10973 17376 10989 17440
rect 11053 17376 11059 17440
rect 10743 17375 11059 17376
rect 15642 17440 15958 17441
rect 15642 17376 15648 17440
rect 15712 17376 15728 17440
rect 15792 17376 15808 17440
rect 15872 17376 15888 17440
rect 15952 17376 15958 17440
rect 15642 17375 15958 17376
rect 20541 17440 20857 17441
rect 20541 17376 20547 17440
rect 20611 17376 20627 17440
rect 20691 17376 20707 17440
rect 20771 17376 20787 17440
rect 20851 17376 20857 17440
rect 20541 17375 20857 17376
rect 3395 16896 3711 16897
rect 3395 16832 3401 16896
rect 3465 16832 3481 16896
rect 3545 16832 3561 16896
rect 3625 16832 3641 16896
rect 3705 16832 3711 16896
rect 3395 16831 3711 16832
rect 8294 16896 8610 16897
rect 8294 16832 8300 16896
rect 8364 16832 8380 16896
rect 8444 16832 8460 16896
rect 8524 16832 8540 16896
rect 8604 16832 8610 16896
rect 8294 16831 8610 16832
rect 13193 16896 13509 16897
rect 13193 16832 13199 16896
rect 13263 16832 13279 16896
rect 13343 16832 13359 16896
rect 13423 16832 13439 16896
rect 13503 16832 13509 16896
rect 13193 16831 13509 16832
rect 18092 16896 18408 16897
rect 18092 16832 18098 16896
rect 18162 16832 18178 16896
rect 18242 16832 18258 16896
rect 18322 16832 18338 16896
rect 18402 16832 18408 16896
rect 18092 16831 18408 16832
rect 20253 16690 20319 16693
rect 21080 16690 21880 16720
rect 20253 16688 21880 16690
rect 20253 16632 20258 16688
rect 20314 16632 21880 16688
rect 20253 16630 21880 16632
rect 20253 16627 20319 16630
rect 21080 16600 21880 16630
rect 5844 16352 6160 16353
rect 5844 16288 5850 16352
rect 5914 16288 5930 16352
rect 5994 16288 6010 16352
rect 6074 16288 6090 16352
rect 6154 16288 6160 16352
rect 5844 16287 6160 16288
rect 10743 16352 11059 16353
rect 10743 16288 10749 16352
rect 10813 16288 10829 16352
rect 10893 16288 10909 16352
rect 10973 16288 10989 16352
rect 11053 16288 11059 16352
rect 10743 16287 11059 16288
rect 15642 16352 15958 16353
rect 15642 16288 15648 16352
rect 15712 16288 15728 16352
rect 15792 16288 15808 16352
rect 15872 16288 15888 16352
rect 15952 16288 15958 16352
rect 15642 16287 15958 16288
rect 20541 16352 20857 16353
rect 20541 16288 20547 16352
rect 20611 16288 20627 16352
rect 20691 16288 20707 16352
rect 20771 16288 20787 16352
rect 20851 16288 20857 16352
rect 20541 16287 20857 16288
rect 3395 15808 3711 15809
rect 3395 15744 3401 15808
rect 3465 15744 3481 15808
rect 3545 15744 3561 15808
rect 3625 15744 3641 15808
rect 3705 15744 3711 15808
rect 3395 15743 3711 15744
rect 8294 15808 8610 15809
rect 8294 15744 8300 15808
rect 8364 15744 8380 15808
rect 8444 15744 8460 15808
rect 8524 15744 8540 15808
rect 8604 15744 8610 15808
rect 8294 15743 8610 15744
rect 13193 15808 13509 15809
rect 13193 15744 13199 15808
rect 13263 15744 13279 15808
rect 13343 15744 13359 15808
rect 13423 15744 13439 15808
rect 13503 15744 13509 15808
rect 13193 15743 13509 15744
rect 18092 15808 18408 15809
rect 18092 15744 18098 15808
rect 18162 15744 18178 15808
rect 18242 15744 18258 15808
rect 18322 15744 18338 15808
rect 18402 15744 18408 15808
rect 18092 15743 18408 15744
rect 5844 15264 6160 15265
rect 5844 15200 5850 15264
rect 5914 15200 5930 15264
rect 5994 15200 6010 15264
rect 6074 15200 6090 15264
rect 6154 15200 6160 15264
rect 5844 15199 6160 15200
rect 10743 15264 11059 15265
rect 10743 15200 10749 15264
rect 10813 15200 10829 15264
rect 10893 15200 10909 15264
rect 10973 15200 10989 15264
rect 11053 15200 11059 15264
rect 10743 15199 11059 15200
rect 15642 15264 15958 15265
rect 15642 15200 15648 15264
rect 15712 15200 15728 15264
rect 15792 15200 15808 15264
rect 15872 15200 15888 15264
rect 15952 15200 15958 15264
rect 15642 15199 15958 15200
rect 20541 15264 20857 15265
rect 20541 15200 20547 15264
rect 20611 15200 20627 15264
rect 20691 15200 20707 15264
rect 20771 15200 20787 15264
rect 20851 15200 20857 15264
rect 20541 15199 20857 15200
rect 19241 15058 19307 15061
rect 21080 15058 21880 15088
rect 19241 15056 21880 15058
rect 19241 15000 19246 15056
rect 19302 15000 21880 15056
rect 19241 14998 21880 15000
rect 19241 14995 19307 14998
rect 21080 14968 21880 14998
rect 3395 14720 3711 14721
rect 3395 14656 3401 14720
rect 3465 14656 3481 14720
rect 3545 14656 3561 14720
rect 3625 14656 3641 14720
rect 3705 14656 3711 14720
rect 3395 14655 3711 14656
rect 8294 14720 8610 14721
rect 8294 14656 8300 14720
rect 8364 14656 8380 14720
rect 8444 14656 8460 14720
rect 8524 14656 8540 14720
rect 8604 14656 8610 14720
rect 8294 14655 8610 14656
rect 13193 14720 13509 14721
rect 13193 14656 13199 14720
rect 13263 14656 13279 14720
rect 13343 14656 13359 14720
rect 13423 14656 13439 14720
rect 13503 14656 13509 14720
rect 13193 14655 13509 14656
rect 18092 14720 18408 14721
rect 18092 14656 18098 14720
rect 18162 14656 18178 14720
rect 18242 14656 18258 14720
rect 18322 14656 18338 14720
rect 18402 14656 18408 14720
rect 18092 14655 18408 14656
rect 5844 14176 6160 14177
rect 5844 14112 5850 14176
rect 5914 14112 5930 14176
rect 5994 14112 6010 14176
rect 6074 14112 6090 14176
rect 6154 14112 6160 14176
rect 5844 14111 6160 14112
rect 10743 14176 11059 14177
rect 10743 14112 10749 14176
rect 10813 14112 10829 14176
rect 10893 14112 10909 14176
rect 10973 14112 10989 14176
rect 11053 14112 11059 14176
rect 10743 14111 11059 14112
rect 15642 14176 15958 14177
rect 15642 14112 15648 14176
rect 15712 14112 15728 14176
rect 15792 14112 15808 14176
rect 15872 14112 15888 14176
rect 15952 14112 15958 14176
rect 15642 14111 15958 14112
rect 20541 14176 20857 14177
rect 20541 14112 20547 14176
rect 20611 14112 20627 14176
rect 20691 14112 20707 14176
rect 20771 14112 20787 14176
rect 20851 14112 20857 14176
rect 20541 14111 20857 14112
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 3395 13632 3711 13633
rect 3395 13568 3401 13632
rect 3465 13568 3481 13632
rect 3545 13568 3561 13632
rect 3625 13568 3641 13632
rect 3705 13568 3711 13632
rect 3395 13567 3711 13568
rect 8294 13632 8610 13633
rect 8294 13568 8300 13632
rect 8364 13568 8380 13632
rect 8444 13568 8460 13632
rect 8524 13568 8540 13632
rect 8604 13568 8610 13632
rect 8294 13567 8610 13568
rect 13193 13632 13509 13633
rect 13193 13568 13199 13632
rect 13263 13568 13279 13632
rect 13343 13568 13359 13632
rect 13423 13568 13439 13632
rect 13503 13568 13509 13632
rect 13193 13567 13509 13568
rect 18092 13632 18408 13633
rect 18092 13568 18098 13632
rect 18162 13568 18178 13632
rect 18242 13568 18258 13632
rect 18322 13568 18338 13632
rect 18402 13568 18408 13632
rect 18092 13567 18408 13568
rect 20161 13426 20227 13429
rect 21080 13426 21880 13456
rect 20161 13424 21880 13426
rect 20161 13368 20166 13424
rect 20222 13368 21880 13424
rect 20161 13366 21880 13368
rect 20161 13363 20227 13366
rect 21080 13336 21880 13366
rect 5844 13088 6160 13089
rect 5844 13024 5850 13088
rect 5914 13024 5930 13088
rect 5994 13024 6010 13088
rect 6074 13024 6090 13088
rect 6154 13024 6160 13088
rect 5844 13023 6160 13024
rect 10743 13088 11059 13089
rect 10743 13024 10749 13088
rect 10813 13024 10829 13088
rect 10893 13024 10909 13088
rect 10973 13024 10989 13088
rect 11053 13024 11059 13088
rect 10743 13023 11059 13024
rect 15642 13088 15958 13089
rect 15642 13024 15648 13088
rect 15712 13024 15728 13088
rect 15792 13024 15808 13088
rect 15872 13024 15888 13088
rect 15952 13024 15958 13088
rect 15642 13023 15958 13024
rect 20541 13088 20857 13089
rect 20541 13024 20547 13088
rect 20611 13024 20627 13088
rect 20691 13024 20707 13088
rect 20771 13024 20787 13088
rect 20851 13024 20857 13088
rect 20541 13023 20857 13024
rect 3395 12544 3711 12545
rect 3395 12480 3401 12544
rect 3465 12480 3481 12544
rect 3545 12480 3561 12544
rect 3625 12480 3641 12544
rect 3705 12480 3711 12544
rect 3395 12479 3711 12480
rect 8294 12544 8610 12545
rect 8294 12480 8300 12544
rect 8364 12480 8380 12544
rect 8444 12480 8460 12544
rect 8524 12480 8540 12544
rect 8604 12480 8610 12544
rect 8294 12479 8610 12480
rect 13193 12544 13509 12545
rect 13193 12480 13199 12544
rect 13263 12480 13279 12544
rect 13343 12480 13359 12544
rect 13423 12480 13439 12544
rect 13503 12480 13509 12544
rect 13193 12479 13509 12480
rect 18092 12544 18408 12545
rect 18092 12480 18098 12544
rect 18162 12480 18178 12544
rect 18242 12480 18258 12544
rect 18322 12480 18338 12544
rect 18402 12480 18408 12544
rect 18092 12479 18408 12480
rect 5844 12000 6160 12001
rect 5844 11936 5850 12000
rect 5914 11936 5930 12000
rect 5994 11936 6010 12000
rect 6074 11936 6090 12000
rect 6154 11936 6160 12000
rect 5844 11935 6160 11936
rect 10743 12000 11059 12001
rect 10743 11936 10749 12000
rect 10813 11936 10829 12000
rect 10893 11936 10909 12000
rect 10973 11936 10989 12000
rect 11053 11936 11059 12000
rect 10743 11935 11059 11936
rect 15642 12000 15958 12001
rect 15642 11936 15648 12000
rect 15712 11936 15728 12000
rect 15792 11936 15808 12000
rect 15872 11936 15888 12000
rect 15952 11936 15958 12000
rect 15642 11935 15958 11936
rect 20541 12000 20857 12001
rect 20541 11936 20547 12000
rect 20611 11936 20627 12000
rect 20691 11936 20707 12000
rect 20771 11936 20787 12000
rect 20851 11936 20857 12000
rect 20541 11935 20857 11936
rect 20161 11794 20227 11797
rect 21080 11794 21880 11824
rect 20161 11792 21880 11794
rect 20161 11736 20166 11792
rect 20222 11736 21880 11792
rect 20161 11734 21880 11736
rect 20161 11731 20227 11734
rect 21080 11704 21880 11734
rect 3395 11456 3711 11457
rect 3395 11392 3401 11456
rect 3465 11392 3481 11456
rect 3545 11392 3561 11456
rect 3625 11392 3641 11456
rect 3705 11392 3711 11456
rect 3395 11391 3711 11392
rect 8294 11456 8610 11457
rect 8294 11392 8300 11456
rect 8364 11392 8380 11456
rect 8444 11392 8460 11456
rect 8524 11392 8540 11456
rect 8604 11392 8610 11456
rect 8294 11391 8610 11392
rect 13193 11456 13509 11457
rect 13193 11392 13199 11456
rect 13263 11392 13279 11456
rect 13343 11392 13359 11456
rect 13423 11392 13439 11456
rect 13503 11392 13509 11456
rect 13193 11391 13509 11392
rect 18092 11456 18408 11457
rect 18092 11392 18098 11456
rect 18162 11392 18178 11456
rect 18242 11392 18258 11456
rect 18322 11392 18338 11456
rect 18402 11392 18408 11456
rect 18092 11391 18408 11392
rect 5844 10912 6160 10913
rect 5844 10848 5850 10912
rect 5914 10848 5930 10912
rect 5994 10848 6010 10912
rect 6074 10848 6090 10912
rect 6154 10848 6160 10912
rect 5844 10847 6160 10848
rect 10743 10912 11059 10913
rect 10743 10848 10749 10912
rect 10813 10848 10829 10912
rect 10893 10848 10909 10912
rect 10973 10848 10989 10912
rect 11053 10848 11059 10912
rect 10743 10847 11059 10848
rect 15642 10912 15958 10913
rect 15642 10848 15648 10912
rect 15712 10848 15728 10912
rect 15792 10848 15808 10912
rect 15872 10848 15888 10912
rect 15952 10848 15958 10912
rect 15642 10847 15958 10848
rect 20541 10912 20857 10913
rect 20541 10848 20547 10912
rect 20611 10848 20627 10912
rect 20691 10848 20707 10912
rect 20771 10848 20787 10912
rect 20851 10848 20857 10912
rect 20541 10847 20857 10848
rect 3395 10368 3711 10369
rect 3395 10304 3401 10368
rect 3465 10304 3481 10368
rect 3545 10304 3561 10368
rect 3625 10304 3641 10368
rect 3705 10304 3711 10368
rect 3395 10303 3711 10304
rect 8294 10368 8610 10369
rect 8294 10304 8300 10368
rect 8364 10304 8380 10368
rect 8444 10304 8460 10368
rect 8524 10304 8540 10368
rect 8604 10304 8610 10368
rect 8294 10303 8610 10304
rect 13193 10368 13509 10369
rect 13193 10304 13199 10368
rect 13263 10304 13279 10368
rect 13343 10304 13359 10368
rect 13423 10304 13439 10368
rect 13503 10304 13509 10368
rect 13193 10303 13509 10304
rect 18092 10368 18408 10369
rect 18092 10304 18098 10368
rect 18162 10304 18178 10368
rect 18242 10304 18258 10368
rect 18322 10304 18338 10368
rect 18402 10304 18408 10368
rect 18092 10303 18408 10304
rect 20161 10162 20227 10165
rect 21080 10162 21880 10192
rect 20161 10160 21880 10162
rect 20161 10104 20166 10160
rect 20222 10104 21880 10160
rect 20161 10102 21880 10104
rect 20161 10099 20227 10102
rect 21080 10072 21880 10102
rect 841 10026 907 10029
rect 798 10024 907 10026
rect 798 9968 846 10024
rect 902 9968 907 10024
rect 798 9963 907 9968
rect 798 9920 858 9963
rect 0 9830 858 9920
rect 0 9800 800 9830
rect 5844 9824 6160 9825
rect 5844 9760 5850 9824
rect 5914 9760 5930 9824
rect 5994 9760 6010 9824
rect 6074 9760 6090 9824
rect 6154 9760 6160 9824
rect 5844 9759 6160 9760
rect 10743 9824 11059 9825
rect 10743 9760 10749 9824
rect 10813 9760 10829 9824
rect 10893 9760 10909 9824
rect 10973 9760 10989 9824
rect 11053 9760 11059 9824
rect 10743 9759 11059 9760
rect 15642 9824 15958 9825
rect 15642 9760 15648 9824
rect 15712 9760 15728 9824
rect 15792 9760 15808 9824
rect 15872 9760 15888 9824
rect 15952 9760 15958 9824
rect 15642 9759 15958 9760
rect 20541 9824 20857 9825
rect 20541 9760 20547 9824
rect 20611 9760 20627 9824
rect 20691 9760 20707 9824
rect 20771 9760 20787 9824
rect 20851 9760 20857 9824
rect 20541 9759 20857 9760
rect 3395 9280 3711 9281
rect 3395 9216 3401 9280
rect 3465 9216 3481 9280
rect 3545 9216 3561 9280
rect 3625 9216 3641 9280
rect 3705 9216 3711 9280
rect 3395 9215 3711 9216
rect 8294 9280 8610 9281
rect 8294 9216 8300 9280
rect 8364 9216 8380 9280
rect 8444 9216 8460 9280
rect 8524 9216 8540 9280
rect 8604 9216 8610 9280
rect 8294 9215 8610 9216
rect 13193 9280 13509 9281
rect 13193 9216 13199 9280
rect 13263 9216 13279 9280
rect 13343 9216 13359 9280
rect 13423 9216 13439 9280
rect 13503 9216 13509 9280
rect 13193 9215 13509 9216
rect 18092 9280 18408 9281
rect 18092 9216 18098 9280
rect 18162 9216 18178 9280
rect 18242 9216 18258 9280
rect 18322 9216 18338 9280
rect 18402 9216 18408 9280
rect 18092 9215 18408 9216
rect 5844 8736 6160 8737
rect 5844 8672 5850 8736
rect 5914 8672 5930 8736
rect 5994 8672 6010 8736
rect 6074 8672 6090 8736
rect 6154 8672 6160 8736
rect 5844 8671 6160 8672
rect 10743 8736 11059 8737
rect 10743 8672 10749 8736
rect 10813 8672 10829 8736
rect 10893 8672 10909 8736
rect 10973 8672 10989 8736
rect 11053 8672 11059 8736
rect 10743 8671 11059 8672
rect 15642 8736 15958 8737
rect 15642 8672 15648 8736
rect 15712 8672 15728 8736
rect 15792 8672 15808 8736
rect 15872 8672 15888 8736
rect 15952 8672 15958 8736
rect 15642 8671 15958 8672
rect 20541 8736 20857 8737
rect 20541 8672 20547 8736
rect 20611 8672 20627 8736
rect 20691 8672 20707 8736
rect 20771 8672 20787 8736
rect 20851 8672 20857 8736
rect 20541 8671 20857 8672
rect 20161 8530 20227 8533
rect 21080 8530 21880 8560
rect 20161 8528 21880 8530
rect 20161 8472 20166 8528
rect 20222 8472 21880 8528
rect 20161 8470 21880 8472
rect 20161 8467 20227 8470
rect 21080 8440 21880 8470
rect 3395 8192 3711 8193
rect 3395 8128 3401 8192
rect 3465 8128 3481 8192
rect 3545 8128 3561 8192
rect 3625 8128 3641 8192
rect 3705 8128 3711 8192
rect 3395 8127 3711 8128
rect 8294 8192 8610 8193
rect 8294 8128 8300 8192
rect 8364 8128 8380 8192
rect 8444 8128 8460 8192
rect 8524 8128 8540 8192
rect 8604 8128 8610 8192
rect 8294 8127 8610 8128
rect 13193 8192 13509 8193
rect 13193 8128 13199 8192
rect 13263 8128 13279 8192
rect 13343 8128 13359 8192
rect 13423 8128 13439 8192
rect 13503 8128 13509 8192
rect 13193 8127 13509 8128
rect 18092 8192 18408 8193
rect 18092 8128 18098 8192
rect 18162 8128 18178 8192
rect 18242 8128 18258 8192
rect 18322 8128 18338 8192
rect 18402 8128 18408 8192
rect 18092 8127 18408 8128
rect 5844 7648 6160 7649
rect 5844 7584 5850 7648
rect 5914 7584 5930 7648
rect 5994 7584 6010 7648
rect 6074 7584 6090 7648
rect 6154 7584 6160 7648
rect 5844 7583 6160 7584
rect 10743 7648 11059 7649
rect 10743 7584 10749 7648
rect 10813 7584 10829 7648
rect 10893 7584 10909 7648
rect 10973 7584 10989 7648
rect 11053 7584 11059 7648
rect 10743 7583 11059 7584
rect 15642 7648 15958 7649
rect 15642 7584 15648 7648
rect 15712 7584 15728 7648
rect 15792 7584 15808 7648
rect 15872 7584 15888 7648
rect 15952 7584 15958 7648
rect 15642 7583 15958 7584
rect 20541 7648 20857 7649
rect 20541 7584 20547 7648
rect 20611 7584 20627 7648
rect 20691 7584 20707 7648
rect 20771 7584 20787 7648
rect 20851 7584 20857 7648
rect 20541 7583 20857 7584
rect 3395 7104 3711 7105
rect 3395 7040 3401 7104
rect 3465 7040 3481 7104
rect 3545 7040 3561 7104
rect 3625 7040 3641 7104
rect 3705 7040 3711 7104
rect 3395 7039 3711 7040
rect 8294 7104 8610 7105
rect 8294 7040 8300 7104
rect 8364 7040 8380 7104
rect 8444 7040 8460 7104
rect 8524 7040 8540 7104
rect 8604 7040 8610 7104
rect 8294 7039 8610 7040
rect 13193 7104 13509 7105
rect 13193 7040 13199 7104
rect 13263 7040 13279 7104
rect 13343 7040 13359 7104
rect 13423 7040 13439 7104
rect 13503 7040 13509 7104
rect 13193 7039 13509 7040
rect 18092 7104 18408 7105
rect 18092 7040 18098 7104
rect 18162 7040 18178 7104
rect 18242 7040 18258 7104
rect 18322 7040 18338 7104
rect 18402 7040 18408 7104
rect 18092 7039 18408 7040
rect 20161 6898 20227 6901
rect 21080 6898 21880 6928
rect 20161 6896 21880 6898
rect 20161 6840 20166 6896
rect 20222 6840 21880 6896
rect 20161 6838 21880 6840
rect 20161 6835 20227 6838
rect 21080 6808 21880 6838
rect 5844 6560 6160 6561
rect 5844 6496 5850 6560
rect 5914 6496 5930 6560
rect 5994 6496 6010 6560
rect 6074 6496 6090 6560
rect 6154 6496 6160 6560
rect 5844 6495 6160 6496
rect 10743 6560 11059 6561
rect 10743 6496 10749 6560
rect 10813 6496 10829 6560
rect 10893 6496 10909 6560
rect 10973 6496 10989 6560
rect 11053 6496 11059 6560
rect 10743 6495 11059 6496
rect 15642 6560 15958 6561
rect 15642 6496 15648 6560
rect 15712 6496 15728 6560
rect 15792 6496 15808 6560
rect 15872 6496 15888 6560
rect 15952 6496 15958 6560
rect 15642 6495 15958 6496
rect 20541 6560 20857 6561
rect 20541 6496 20547 6560
rect 20611 6496 20627 6560
rect 20691 6496 20707 6560
rect 20771 6496 20787 6560
rect 20851 6496 20857 6560
rect 20541 6495 20857 6496
rect 4889 6218 4955 6221
rect 2454 6216 4955 6218
rect 2454 6160 4894 6216
rect 4950 6160 4955 6216
rect 2454 6158 4955 6160
rect 0 6082 800 6112
rect 2454 6082 2514 6158
rect 4889 6155 4955 6158
rect 0 6022 2514 6082
rect 0 5992 800 6022
rect 3395 6016 3711 6017
rect 3395 5952 3401 6016
rect 3465 5952 3481 6016
rect 3545 5952 3561 6016
rect 3625 5952 3641 6016
rect 3705 5952 3711 6016
rect 3395 5951 3711 5952
rect 8294 6016 8610 6017
rect 8294 5952 8300 6016
rect 8364 5952 8380 6016
rect 8444 5952 8460 6016
rect 8524 5952 8540 6016
rect 8604 5952 8610 6016
rect 8294 5951 8610 5952
rect 13193 6016 13509 6017
rect 13193 5952 13199 6016
rect 13263 5952 13279 6016
rect 13343 5952 13359 6016
rect 13423 5952 13439 6016
rect 13503 5952 13509 6016
rect 13193 5951 13509 5952
rect 18092 6016 18408 6017
rect 18092 5952 18098 6016
rect 18162 5952 18178 6016
rect 18242 5952 18258 6016
rect 18322 5952 18338 6016
rect 18402 5952 18408 6016
rect 18092 5951 18408 5952
rect 5844 5472 6160 5473
rect 5844 5408 5850 5472
rect 5914 5408 5930 5472
rect 5994 5408 6010 5472
rect 6074 5408 6090 5472
rect 6154 5408 6160 5472
rect 5844 5407 6160 5408
rect 10743 5472 11059 5473
rect 10743 5408 10749 5472
rect 10813 5408 10829 5472
rect 10893 5408 10909 5472
rect 10973 5408 10989 5472
rect 11053 5408 11059 5472
rect 10743 5407 11059 5408
rect 15642 5472 15958 5473
rect 15642 5408 15648 5472
rect 15712 5408 15728 5472
rect 15792 5408 15808 5472
rect 15872 5408 15888 5472
rect 15952 5408 15958 5472
rect 15642 5407 15958 5408
rect 20541 5472 20857 5473
rect 20541 5408 20547 5472
rect 20611 5408 20627 5472
rect 20691 5408 20707 5472
rect 20771 5408 20787 5472
rect 20851 5408 20857 5472
rect 20541 5407 20857 5408
rect 20253 5266 20319 5269
rect 21080 5266 21880 5296
rect 20253 5264 21880 5266
rect 20253 5208 20258 5264
rect 20314 5208 21880 5264
rect 20253 5206 21880 5208
rect 20253 5203 20319 5206
rect 21080 5176 21880 5206
rect 3395 4928 3711 4929
rect 3395 4864 3401 4928
rect 3465 4864 3481 4928
rect 3545 4864 3561 4928
rect 3625 4864 3641 4928
rect 3705 4864 3711 4928
rect 3395 4863 3711 4864
rect 8294 4928 8610 4929
rect 8294 4864 8300 4928
rect 8364 4864 8380 4928
rect 8444 4864 8460 4928
rect 8524 4864 8540 4928
rect 8604 4864 8610 4928
rect 8294 4863 8610 4864
rect 13193 4928 13509 4929
rect 13193 4864 13199 4928
rect 13263 4864 13279 4928
rect 13343 4864 13359 4928
rect 13423 4864 13439 4928
rect 13503 4864 13509 4928
rect 13193 4863 13509 4864
rect 18092 4928 18408 4929
rect 18092 4864 18098 4928
rect 18162 4864 18178 4928
rect 18242 4864 18258 4928
rect 18322 4864 18338 4928
rect 18402 4864 18408 4928
rect 18092 4863 18408 4864
rect 5844 4384 6160 4385
rect 5844 4320 5850 4384
rect 5914 4320 5930 4384
rect 5994 4320 6010 4384
rect 6074 4320 6090 4384
rect 6154 4320 6160 4384
rect 5844 4319 6160 4320
rect 10743 4384 11059 4385
rect 10743 4320 10749 4384
rect 10813 4320 10829 4384
rect 10893 4320 10909 4384
rect 10973 4320 10989 4384
rect 11053 4320 11059 4384
rect 10743 4319 11059 4320
rect 15642 4384 15958 4385
rect 15642 4320 15648 4384
rect 15712 4320 15728 4384
rect 15792 4320 15808 4384
rect 15872 4320 15888 4384
rect 15952 4320 15958 4384
rect 15642 4319 15958 4320
rect 20541 4384 20857 4385
rect 20541 4320 20547 4384
rect 20611 4320 20627 4384
rect 20691 4320 20707 4384
rect 20771 4320 20787 4384
rect 20851 4320 20857 4384
rect 20541 4319 20857 4320
rect 3395 3840 3711 3841
rect 3395 3776 3401 3840
rect 3465 3776 3481 3840
rect 3545 3776 3561 3840
rect 3625 3776 3641 3840
rect 3705 3776 3711 3840
rect 3395 3775 3711 3776
rect 8294 3840 8610 3841
rect 8294 3776 8300 3840
rect 8364 3776 8380 3840
rect 8444 3776 8460 3840
rect 8524 3776 8540 3840
rect 8604 3776 8610 3840
rect 8294 3775 8610 3776
rect 13193 3840 13509 3841
rect 13193 3776 13199 3840
rect 13263 3776 13279 3840
rect 13343 3776 13359 3840
rect 13423 3776 13439 3840
rect 13503 3776 13509 3840
rect 13193 3775 13509 3776
rect 18092 3840 18408 3841
rect 18092 3776 18098 3840
rect 18162 3776 18178 3840
rect 18242 3776 18258 3840
rect 18322 3776 18338 3840
rect 18402 3776 18408 3840
rect 18092 3775 18408 3776
rect 20253 3634 20319 3637
rect 21080 3634 21880 3664
rect 20253 3632 21880 3634
rect 20253 3576 20258 3632
rect 20314 3576 21880 3632
rect 20253 3574 21880 3576
rect 20253 3571 20319 3574
rect 21080 3544 21880 3574
rect 5844 3296 6160 3297
rect 5844 3232 5850 3296
rect 5914 3232 5930 3296
rect 5994 3232 6010 3296
rect 6074 3232 6090 3296
rect 6154 3232 6160 3296
rect 5844 3231 6160 3232
rect 10743 3296 11059 3297
rect 10743 3232 10749 3296
rect 10813 3232 10829 3296
rect 10893 3232 10909 3296
rect 10973 3232 10989 3296
rect 11053 3232 11059 3296
rect 10743 3231 11059 3232
rect 15642 3296 15958 3297
rect 15642 3232 15648 3296
rect 15712 3232 15728 3296
rect 15792 3232 15808 3296
rect 15872 3232 15888 3296
rect 15952 3232 15958 3296
rect 15642 3231 15958 3232
rect 20541 3296 20857 3297
rect 20541 3232 20547 3296
rect 20611 3232 20627 3296
rect 20691 3232 20707 3296
rect 20771 3232 20787 3296
rect 20851 3232 20857 3296
rect 20541 3231 20857 3232
rect 3395 2752 3711 2753
rect 3395 2688 3401 2752
rect 3465 2688 3481 2752
rect 3545 2688 3561 2752
rect 3625 2688 3641 2752
rect 3705 2688 3711 2752
rect 3395 2687 3711 2688
rect 8294 2752 8610 2753
rect 8294 2688 8300 2752
rect 8364 2688 8380 2752
rect 8444 2688 8460 2752
rect 8524 2688 8540 2752
rect 8604 2688 8610 2752
rect 8294 2687 8610 2688
rect 13193 2752 13509 2753
rect 13193 2688 13199 2752
rect 13263 2688 13279 2752
rect 13343 2688 13359 2752
rect 13423 2688 13439 2752
rect 13503 2688 13509 2752
rect 13193 2687 13509 2688
rect 18092 2752 18408 2753
rect 18092 2688 18098 2752
rect 18162 2688 18178 2752
rect 18242 2688 18258 2752
rect 18322 2688 18338 2752
rect 18402 2688 18408 2752
rect 18092 2687 18408 2688
rect 0 2274 800 2304
rect 1485 2274 1551 2277
rect 0 2272 1551 2274
rect 0 2216 1490 2272
rect 1546 2216 1551 2272
rect 0 2214 1551 2216
rect 0 2184 800 2214
rect 1485 2211 1551 2214
rect 5844 2208 6160 2209
rect 5844 2144 5850 2208
rect 5914 2144 5930 2208
rect 5994 2144 6010 2208
rect 6074 2144 6090 2208
rect 6154 2144 6160 2208
rect 5844 2143 6160 2144
rect 10743 2208 11059 2209
rect 10743 2144 10749 2208
rect 10813 2144 10829 2208
rect 10893 2144 10909 2208
rect 10973 2144 10989 2208
rect 11053 2144 11059 2208
rect 10743 2143 11059 2144
rect 15642 2208 15958 2209
rect 15642 2144 15648 2208
rect 15712 2144 15728 2208
rect 15792 2144 15808 2208
rect 15872 2144 15888 2208
rect 15952 2144 15958 2208
rect 15642 2143 15958 2144
rect 20541 2208 20857 2209
rect 20541 2144 20547 2208
rect 20611 2144 20627 2208
rect 20691 2144 20707 2208
rect 20771 2144 20787 2208
rect 20851 2144 20857 2208
rect 20541 2143 20857 2144
rect 20161 2002 20227 2005
rect 21080 2002 21880 2032
rect 20161 2000 21880 2002
rect 20161 1944 20166 2000
rect 20222 1944 21880 2000
rect 20161 1942 21880 1944
rect 20161 1939 20227 1942
rect 21080 1912 21880 1942
<< via3 >>
rect 5850 21788 5914 21792
rect 5850 21732 5854 21788
rect 5854 21732 5910 21788
rect 5910 21732 5914 21788
rect 5850 21728 5914 21732
rect 5930 21788 5994 21792
rect 5930 21732 5934 21788
rect 5934 21732 5990 21788
rect 5990 21732 5994 21788
rect 5930 21728 5994 21732
rect 6010 21788 6074 21792
rect 6010 21732 6014 21788
rect 6014 21732 6070 21788
rect 6070 21732 6074 21788
rect 6010 21728 6074 21732
rect 6090 21788 6154 21792
rect 6090 21732 6094 21788
rect 6094 21732 6150 21788
rect 6150 21732 6154 21788
rect 6090 21728 6154 21732
rect 10749 21788 10813 21792
rect 10749 21732 10753 21788
rect 10753 21732 10809 21788
rect 10809 21732 10813 21788
rect 10749 21728 10813 21732
rect 10829 21788 10893 21792
rect 10829 21732 10833 21788
rect 10833 21732 10889 21788
rect 10889 21732 10893 21788
rect 10829 21728 10893 21732
rect 10909 21788 10973 21792
rect 10909 21732 10913 21788
rect 10913 21732 10969 21788
rect 10969 21732 10973 21788
rect 10909 21728 10973 21732
rect 10989 21788 11053 21792
rect 10989 21732 10993 21788
rect 10993 21732 11049 21788
rect 11049 21732 11053 21788
rect 10989 21728 11053 21732
rect 15648 21788 15712 21792
rect 15648 21732 15652 21788
rect 15652 21732 15708 21788
rect 15708 21732 15712 21788
rect 15648 21728 15712 21732
rect 15728 21788 15792 21792
rect 15728 21732 15732 21788
rect 15732 21732 15788 21788
rect 15788 21732 15792 21788
rect 15728 21728 15792 21732
rect 15808 21788 15872 21792
rect 15808 21732 15812 21788
rect 15812 21732 15868 21788
rect 15868 21732 15872 21788
rect 15808 21728 15872 21732
rect 15888 21788 15952 21792
rect 15888 21732 15892 21788
rect 15892 21732 15948 21788
rect 15948 21732 15952 21788
rect 15888 21728 15952 21732
rect 20547 21788 20611 21792
rect 20547 21732 20551 21788
rect 20551 21732 20607 21788
rect 20607 21732 20611 21788
rect 20547 21728 20611 21732
rect 20627 21788 20691 21792
rect 20627 21732 20631 21788
rect 20631 21732 20687 21788
rect 20687 21732 20691 21788
rect 20627 21728 20691 21732
rect 20707 21788 20771 21792
rect 20707 21732 20711 21788
rect 20711 21732 20767 21788
rect 20767 21732 20771 21788
rect 20707 21728 20771 21732
rect 20787 21788 20851 21792
rect 20787 21732 20791 21788
rect 20791 21732 20847 21788
rect 20847 21732 20851 21788
rect 20787 21728 20851 21732
rect 3401 21244 3465 21248
rect 3401 21188 3405 21244
rect 3405 21188 3461 21244
rect 3461 21188 3465 21244
rect 3401 21184 3465 21188
rect 3481 21244 3545 21248
rect 3481 21188 3485 21244
rect 3485 21188 3541 21244
rect 3541 21188 3545 21244
rect 3481 21184 3545 21188
rect 3561 21244 3625 21248
rect 3561 21188 3565 21244
rect 3565 21188 3621 21244
rect 3621 21188 3625 21244
rect 3561 21184 3625 21188
rect 3641 21244 3705 21248
rect 3641 21188 3645 21244
rect 3645 21188 3701 21244
rect 3701 21188 3705 21244
rect 3641 21184 3705 21188
rect 8300 21244 8364 21248
rect 8300 21188 8304 21244
rect 8304 21188 8360 21244
rect 8360 21188 8364 21244
rect 8300 21184 8364 21188
rect 8380 21244 8444 21248
rect 8380 21188 8384 21244
rect 8384 21188 8440 21244
rect 8440 21188 8444 21244
rect 8380 21184 8444 21188
rect 8460 21244 8524 21248
rect 8460 21188 8464 21244
rect 8464 21188 8520 21244
rect 8520 21188 8524 21244
rect 8460 21184 8524 21188
rect 8540 21244 8604 21248
rect 8540 21188 8544 21244
rect 8544 21188 8600 21244
rect 8600 21188 8604 21244
rect 8540 21184 8604 21188
rect 13199 21244 13263 21248
rect 13199 21188 13203 21244
rect 13203 21188 13259 21244
rect 13259 21188 13263 21244
rect 13199 21184 13263 21188
rect 13279 21244 13343 21248
rect 13279 21188 13283 21244
rect 13283 21188 13339 21244
rect 13339 21188 13343 21244
rect 13279 21184 13343 21188
rect 13359 21244 13423 21248
rect 13359 21188 13363 21244
rect 13363 21188 13419 21244
rect 13419 21188 13423 21244
rect 13359 21184 13423 21188
rect 13439 21244 13503 21248
rect 13439 21188 13443 21244
rect 13443 21188 13499 21244
rect 13499 21188 13503 21244
rect 13439 21184 13503 21188
rect 18098 21244 18162 21248
rect 18098 21188 18102 21244
rect 18102 21188 18158 21244
rect 18158 21188 18162 21244
rect 18098 21184 18162 21188
rect 18178 21244 18242 21248
rect 18178 21188 18182 21244
rect 18182 21188 18238 21244
rect 18238 21188 18242 21244
rect 18178 21184 18242 21188
rect 18258 21244 18322 21248
rect 18258 21188 18262 21244
rect 18262 21188 18318 21244
rect 18318 21188 18322 21244
rect 18258 21184 18322 21188
rect 18338 21244 18402 21248
rect 18338 21188 18342 21244
rect 18342 21188 18398 21244
rect 18398 21188 18402 21244
rect 18338 21184 18402 21188
rect 5850 20700 5914 20704
rect 5850 20644 5854 20700
rect 5854 20644 5910 20700
rect 5910 20644 5914 20700
rect 5850 20640 5914 20644
rect 5930 20700 5994 20704
rect 5930 20644 5934 20700
rect 5934 20644 5990 20700
rect 5990 20644 5994 20700
rect 5930 20640 5994 20644
rect 6010 20700 6074 20704
rect 6010 20644 6014 20700
rect 6014 20644 6070 20700
rect 6070 20644 6074 20700
rect 6010 20640 6074 20644
rect 6090 20700 6154 20704
rect 6090 20644 6094 20700
rect 6094 20644 6150 20700
rect 6150 20644 6154 20700
rect 6090 20640 6154 20644
rect 10749 20700 10813 20704
rect 10749 20644 10753 20700
rect 10753 20644 10809 20700
rect 10809 20644 10813 20700
rect 10749 20640 10813 20644
rect 10829 20700 10893 20704
rect 10829 20644 10833 20700
rect 10833 20644 10889 20700
rect 10889 20644 10893 20700
rect 10829 20640 10893 20644
rect 10909 20700 10973 20704
rect 10909 20644 10913 20700
rect 10913 20644 10969 20700
rect 10969 20644 10973 20700
rect 10909 20640 10973 20644
rect 10989 20700 11053 20704
rect 10989 20644 10993 20700
rect 10993 20644 11049 20700
rect 11049 20644 11053 20700
rect 10989 20640 11053 20644
rect 15648 20700 15712 20704
rect 15648 20644 15652 20700
rect 15652 20644 15708 20700
rect 15708 20644 15712 20700
rect 15648 20640 15712 20644
rect 15728 20700 15792 20704
rect 15728 20644 15732 20700
rect 15732 20644 15788 20700
rect 15788 20644 15792 20700
rect 15728 20640 15792 20644
rect 15808 20700 15872 20704
rect 15808 20644 15812 20700
rect 15812 20644 15868 20700
rect 15868 20644 15872 20700
rect 15808 20640 15872 20644
rect 15888 20700 15952 20704
rect 15888 20644 15892 20700
rect 15892 20644 15948 20700
rect 15948 20644 15952 20700
rect 15888 20640 15952 20644
rect 20547 20700 20611 20704
rect 20547 20644 20551 20700
rect 20551 20644 20607 20700
rect 20607 20644 20611 20700
rect 20547 20640 20611 20644
rect 20627 20700 20691 20704
rect 20627 20644 20631 20700
rect 20631 20644 20687 20700
rect 20687 20644 20691 20700
rect 20627 20640 20691 20644
rect 20707 20700 20771 20704
rect 20707 20644 20711 20700
rect 20711 20644 20767 20700
rect 20767 20644 20771 20700
rect 20707 20640 20771 20644
rect 20787 20700 20851 20704
rect 20787 20644 20791 20700
rect 20791 20644 20847 20700
rect 20847 20644 20851 20700
rect 20787 20640 20851 20644
rect 3401 20156 3465 20160
rect 3401 20100 3405 20156
rect 3405 20100 3461 20156
rect 3461 20100 3465 20156
rect 3401 20096 3465 20100
rect 3481 20156 3545 20160
rect 3481 20100 3485 20156
rect 3485 20100 3541 20156
rect 3541 20100 3545 20156
rect 3481 20096 3545 20100
rect 3561 20156 3625 20160
rect 3561 20100 3565 20156
rect 3565 20100 3621 20156
rect 3621 20100 3625 20156
rect 3561 20096 3625 20100
rect 3641 20156 3705 20160
rect 3641 20100 3645 20156
rect 3645 20100 3701 20156
rect 3701 20100 3705 20156
rect 3641 20096 3705 20100
rect 8300 20156 8364 20160
rect 8300 20100 8304 20156
rect 8304 20100 8360 20156
rect 8360 20100 8364 20156
rect 8300 20096 8364 20100
rect 8380 20156 8444 20160
rect 8380 20100 8384 20156
rect 8384 20100 8440 20156
rect 8440 20100 8444 20156
rect 8380 20096 8444 20100
rect 8460 20156 8524 20160
rect 8460 20100 8464 20156
rect 8464 20100 8520 20156
rect 8520 20100 8524 20156
rect 8460 20096 8524 20100
rect 8540 20156 8604 20160
rect 8540 20100 8544 20156
rect 8544 20100 8600 20156
rect 8600 20100 8604 20156
rect 8540 20096 8604 20100
rect 13199 20156 13263 20160
rect 13199 20100 13203 20156
rect 13203 20100 13259 20156
rect 13259 20100 13263 20156
rect 13199 20096 13263 20100
rect 13279 20156 13343 20160
rect 13279 20100 13283 20156
rect 13283 20100 13339 20156
rect 13339 20100 13343 20156
rect 13279 20096 13343 20100
rect 13359 20156 13423 20160
rect 13359 20100 13363 20156
rect 13363 20100 13419 20156
rect 13419 20100 13423 20156
rect 13359 20096 13423 20100
rect 13439 20156 13503 20160
rect 13439 20100 13443 20156
rect 13443 20100 13499 20156
rect 13499 20100 13503 20156
rect 13439 20096 13503 20100
rect 18098 20156 18162 20160
rect 18098 20100 18102 20156
rect 18102 20100 18158 20156
rect 18158 20100 18162 20156
rect 18098 20096 18162 20100
rect 18178 20156 18242 20160
rect 18178 20100 18182 20156
rect 18182 20100 18238 20156
rect 18238 20100 18242 20156
rect 18178 20096 18242 20100
rect 18258 20156 18322 20160
rect 18258 20100 18262 20156
rect 18262 20100 18318 20156
rect 18318 20100 18322 20156
rect 18258 20096 18322 20100
rect 18338 20156 18402 20160
rect 18338 20100 18342 20156
rect 18342 20100 18398 20156
rect 18398 20100 18402 20156
rect 18338 20096 18402 20100
rect 5850 19612 5914 19616
rect 5850 19556 5854 19612
rect 5854 19556 5910 19612
rect 5910 19556 5914 19612
rect 5850 19552 5914 19556
rect 5930 19612 5994 19616
rect 5930 19556 5934 19612
rect 5934 19556 5990 19612
rect 5990 19556 5994 19612
rect 5930 19552 5994 19556
rect 6010 19612 6074 19616
rect 6010 19556 6014 19612
rect 6014 19556 6070 19612
rect 6070 19556 6074 19612
rect 6010 19552 6074 19556
rect 6090 19612 6154 19616
rect 6090 19556 6094 19612
rect 6094 19556 6150 19612
rect 6150 19556 6154 19612
rect 6090 19552 6154 19556
rect 10749 19612 10813 19616
rect 10749 19556 10753 19612
rect 10753 19556 10809 19612
rect 10809 19556 10813 19612
rect 10749 19552 10813 19556
rect 10829 19612 10893 19616
rect 10829 19556 10833 19612
rect 10833 19556 10889 19612
rect 10889 19556 10893 19612
rect 10829 19552 10893 19556
rect 10909 19612 10973 19616
rect 10909 19556 10913 19612
rect 10913 19556 10969 19612
rect 10969 19556 10973 19612
rect 10909 19552 10973 19556
rect 10989 19612 11053 19616
rect 10989 19556 10993 19612
rect 10993 19556 11049 19612
rect 11049 19556 11053 19612
rect 10989 19552 11053 19556
rect 15648 19612 15712 19616
rect 15648 19556 15652 19612
rect 15652 19556 15708 19612
rect 15708 19556 15712 19612
rect 15648 19552 15712 19556
rect 15728 19612 15792 19616
rect 15728 19556 15732 19612
rect 15732 19556 15788 19612
rect 15788 19556 15792 19612
rect 15728 19552 15792 19556
rect 15808 19612 15872 19616
rect 15808 19556 15812 19612
rect 15812 19556 15868 19612
rect 15868 19556 15872 19612
rect 15808 19552 15872 19556
rect 15888 19612 15952 19616
rect 15888 19556 15892 19612
rect 15892 19556 15948 19612
rect 15948 19556 15952 19612
rect 15888 19552 15952 19556
rect 20547 19612 20611 19616
rect 20547 19556 20551 19612
rect 20551 19556 20607 19612
rect 20607 19556 20611 19612
rect 20547 19552 20611 19556
rect 20627 19612 20691 19616
rect 20627 19556 20631 19612
rect 20631 19556 20687 19612
rect 20687 19556 20691 19612
rect 20627 19552 20691 19556
rect 20707 19612 20771 19616
rect 20707 19556 20711 19612
rect 20711 19556 20767 19612
rect 20767 19556 20771 19612
rect 20707 19552 20771 19556
rect 20787 19612 20851 19616
rect 20787 19556 20791 19612
rect 20791 19556 20847 19612
rect 20847 19556 20851 19612
rect 20787 19552 20851 19556
rect 3401 19068 3465 19072
rect 3401 19012 3405 19068
rect 3405 19012 3461 19068
rect 3461 19012 3465 19068
rect 3401 19008 3465 19012
rect 3481 19068 3545 19072
rect 3481 19012 3485 19068
rect 3485 19012 3541 19068
rect 3541 19012 3545 19068
rect 3481 19008 3545 19012
rect 3561 19068 3625 19072
rect 3561 19012 3565 19068
rect 3565 19012 3621 19068
rect 3621 19012 3625 19068
rect 3561 19008 3625 19012
rect 3641 19068 3705 19072
rect 3641 19012 3645 19068
rect 3645 19012 3701 19068
rect 3701 19012 3705 19068
rect 3641 19008 3705 19012
rect 8300 19068 8364 19072
rect 8300 19012 8304 19068
rect 8304 19012 8360 19068
rect 8360 19012 8364 19068
rect 8300 19008 8364 19012
rect 8380 19068 8444 19072
rect 8380 19012 8384 19068
rect 8384 19012 8440 19068
rect 8440 19012 8444 19068
rect 8380 19008 8444 19012
rect 8460 19068 8524 19072
rect 8460 19012 8464 19068
rect 8464 19012 8520 19068
rect 8520 19012 8524 19068
rect 8460 19008 8524 19012
rect 8540 19068 8604 19072
rect 8540 19012 8544 19068
rect 8544 19012 8600 19068
rect 8600 19012 8604 19068
rect 8540 19008 8604 19012
rect 13199 19068 13263 19072
rect 13199 19012 13203 19068
rect 13203 19012 13259 19068
rect 13259 19012 13263 19068
rect 13199 19008 13263 19012
rect 13279 19068 13343 19072
rect 13279 19012 13283 19068
rect 13283 19012 13339 19068
rect 13339 19012 13343 19068
rect 13279 19008 13343 19012
rect 13359 19068 13423 19072
rect 13359 19012 13363 19068
rect 13363 19012 13419 19068
rect 13419 19012 13423 19068
rect 13359 19008 13423 19012
rect 13439 19068 13503 19072
rect 13439 19012 13443 19068
rect 13443 19012 13499 19068
rect 13499 19012 13503 19068
rect 13439 19008 13503 19012
rect 18098 19068 18162 19072
rect 18098 19012 18102 19068
rect 18102 19012 18158 19068
rect 18158 19012 18162 19068
rect 18098 19008 18162 19012
rect 18178 19068 18242 19072
rect 18178 19012 18182 19068
rect 18182 19012 18238 19068
rect 18238 19012 18242 19068
rect 18178 19008 18242 19012
rect 18258 19068 18322 19072
rect 18258 19012 18262 19068
rect 18262 19012 18318 19068
rect 18318 19012 18322 19068
rect 18258 19008 18322 19012
rect 18338 19068 18402 19072
rect 18338 19012 18342 19068
rect 18342 19012 18398 19068
rect 18398 19012 18402 19068
rect 18338 19008 18402 19012
rect 5850 18524 5914 18528
rect 5850 18468 5854 18524
rect 5854 18468 5910 18524
rect 5910 18468 5914 18524
rect 5850 18464 5914 18468
rect 5930 18524 5994 18528
rect 5930 18468 5934 18524
rect 5934 18468 5990 18524
rect 5990 18468 5994 18524
rect 5930 18464 5994 18468
rect 6010 18524 6074 18528
rect 6010 18468 6014 18524
rect 6014 18468 6070 18524
rect 6070 18468 6074 18524
rect 6010 18464 6074 18468
rect 6090 18524 6154 18528
rect 6090 18468 6094 18524
rect 6094 18468 6150 18524
rect 6150 18468 6154 18524
rect 6090 18464 6154 18468
rect 10749 18524 10813 18528
rect 10749 18468 10753 18524
rect 10753 18468 10809 18524
rect 10809 18468 10813 18524
rect 10749 18464 10813 18468
rect 10829 18524 10893 18528
rect 10829 18468 10833 18524
rect 10833 18468 10889 18524
rect 10889 18468 10893 18524
rect 10829 18464 10893 18468
rect 10909 18524 10973 18528
rect 10909 18468 10913 18524
rect 10913 18468 10969 18524
rect 10969 18468 10973 18524
rect 10909 18464 10973 18468
rect 10989 18524 11053 18528
rect 10989 18468 10993 18524
rect 10993 18468 11049 18524
rect 11049 18468 11053 18524
rect 10989 18464 11053 18468
rect 15648 18524 15712 18528
rect 15648 18468 15652 18524
rect 15652 18468 15708 18524
rect 15708 18468 15712 18524
rect 15648 18464 15712 18468
rect 15728 18524 15792 18528
rect 15728 18468 15732 18524
rect 15732 18468 15788 18524
rect 15788 18468 15792 18524
rect 15728 18464 15792 18468
rect 15808 18524 15872 18528
rect 15808 18468 15812 18524
rect 15812 18468 15868 18524
rect 15868 18468 15872 18524
rect 15808 18464 15872 18468
rect 15888 18524 15952 18528
rect 15888 18468 15892 18524
rect 15892 18468 15948 18524
rect 15948 18468 15952 18524
rect 15888 18464 15952 18468
rect 20547 18524 20611 18528
rect 20547 18468 20551 18524
rect 20551 18468 20607 18524
rect 20607 18468 20611 18524
rect 20547 18464 20611 18468
rect 20627 18524 20691 18528
rect 20627 18468 20631 18524
rect 20631 18468 20687 18524
rect 20687 18468 20691 18524
rect 20627 18464 20691 18468
rect 20707 18524 20771 18528
rect 20707 18468 20711 18524
rect 20711 18468 20767 18524
rect 20767 18468 20771 18524
rect 20707 18464 20771 18468
rect 20787 18524 20851 18528
rect 20787 18468 20791 18524
rect 20791 18468 20847 18524
rect 20847 18468 20851 18524
rect 20787 18464 20851 18468
rect 3401 17980 3465 17984
rect 3401 17924 3405 17980
rect 3405 17924 3461 17980
rect 3461 17924 3465 17980
rect 3401 17920 3465 17924
rect 3481 17980 3545 17984
rect 3481 17924 3485 17980
rect 3485 17924 3541 17980
rect 3541 17924 3545 17980
rect 3481 17920 3545 17924
rect 3561 17980 3625 17984
rect 3561 17924 3565 17980
rect 3565 17924 3621 17980
rect 3621 17924 3625 17980
rect 3561 17920 3625 17924
rect 3641 17980 3705 17984
rect 3641 17924 3645 17980
rect 3645 17924 3701 17980
rect 3701 17924 3705 17980
rect 3641 17920 3705 17924
rect 8300 17980 8364 17984
rect 8300 17924 8304 17980
rect 8304 17924 8360 17980
rect 8360 17924 8364 17980
rect 8300 17920 8364 17924
rect 8380 17980 8444 17984
rect 8380 17924 8384 17980
rect 8384 17924 8440 17980
rect 8440 17924 8444 17980
rect 8380 17920 8444 17924
rect 8460 17980 8524 17984
rect 8460 17924 8464 17980
rect 8464 17924 8520 17980
rect 8520 17924 8524 17980
rect 8460 17920 8524 17924
rect 8540 17980 8604 17984
rect 8540 17924 8544 17980
rect 8544 17924 8600 17980
rect 8600 17924 8604 17980
rect 8540 17920 8604 17924
rect 13199 17980 13263 17984
rect 13199 17924 13203 17980
rect 13203 17924 13259 17980
rect 13259 17924 13263 17980
rect 13199 17920 13263 17924
rect 13279 17980 13343 17984
rect 13279 17924 13283 17980
rect 13283 17924 13339 17980
rect 13339 17924 13343 17980
rect 13279 17920 13343 17924
rect 13359 17980 13423 17984
rect 13359 17924 13363 17980
rect 13363 17924 13419 17980
rect 13419 17924 13423 17980
rect 13359 17920 13423 17924
rect 13439 17980 13503 17984
rect 13439 17924 13443 17980
rect 13443 17924 13499 17980
rect 13499 17924 13503 17980
rect 13439 17920 13503 17924
rect 18098 17980 18162 17984
rect 18098 17924 18102 17980
rect 18102 17924 18158 17980
rect 18158 17924 18162 17980
rect 18098 17920 18162 17924
rect 18178 17980 18242 17984
rect 18178 17924 18182 17980
rect 18182 17924 18238 17980
rect 18238 17924 18242 17980
rect 18178 17920 18242 17924
rect 18258 17980 18322 17984
rect 18258 17924 18262 17980
rect 18262 17924 18318 17980
rect 18318 17924 18322 17980
rect 18258 17920 18322 17924
rect 18338 17980 18402 17984
rect 18338 17924 18342 17980
rect 18342 17924 18398 17980
rect 18398 17924 18402 17980
rect 18338 17920 18402 17924
rect 5850 17436 5914 17440
rect 5850 17380 5854 17436
rect 5854 17380 5910 17436
rect 5910 17380 5914 17436
rect 5850 17376 5914 17380
rect 5930 17436 5994 17440
rect 5930 17380 5934 17436
rect 5934 17380 5990 17436
rect 5990 17380 5994 17436
rect 5930 17376 5994 17380
rect 6010 17436 6074 17440
rect 6010 17380 6014 17436
rect 6014 17380 6070 17436
rect 6070 17380 6074 17436
rect 6010 17376 6074 17380
rect 6090 17436 6154 17440
rect 6090 17380 6094 17436
rect 6094 17380 6150 17436
rect 6150 17380 6154 17436
rect 6090 17376 6154 17380
rect 10749 17436 10813 17440
rect 10749 17380 10753 17436
rect 10753 17380 10809 17436
rect 10809 17380 10813 17436
rect 10749 17376 10813 17380
rect 10829 17436 10893 17440
rect 10829 17380 10833 17436
rect 10833 17380 10889 17436
rect 10889 17380 10893 17436
rect 10829 17376 10893 17380
rect 10909 17436 10973 17440
rect 10909 17380 10913 17436
rect 10913 17380 10969 17436
rect 10969 17380 10973 17436
rect 10909 17376 10973 17380
rect 10989 17436 11053 17440
rect 10989 17380 10993 17436
rect 10993 17380 11049 17436
rect 11049 17380 11053 17436
rect 10989 17376 11053 17380
rect 15648 17436 15712 17440
rect 15648 17380 15652 17436
rect 15652 17380 15708 17436
rect 15708 17380 15712 17436
rect 15648 17376 15712 17380
rect 15728 17436 15792 17440
rect 15728 17380 15732 17436
rect 15732 17380 15788 17436
rect 15788 17380 15792 17436
rect 15728 17376 15792 17380
rect 15808 17436 15872 17440
rect 15808 17380 15812 17436
rect 15812 17380 15868 17436
rect 15868 17380 15872 17436
rect 15808 17376 15872 17380
rect 15888 17436 15952 17440
rect 15888 17380 15892 17436
rect 15892 17380 15948 17436
rect 15948 17380 15952 17436
rect 15888 17376 15952 17380
rect 20547 17436 20611 17440
rect 20547 17380 20551 17436
rect 20551 17380 20607 17436
rect 20607 17380 20611 17436
rect 20547 17376 20611 17380
rect 20627 17436 20691 17440
rect 20627 17380 20631 17436
rect 20631 17380 20687 17436
rect 20687 17380 20691 17436
rect 20627 17376 20691 17380
rect 20707 17436 20771 17440
rect 20707 17380 20711 17436
rect 20711 17380 20767 17436
rect 20767 17380 20771 17436
rect 20707 17376 20771 17380
rect 20787 17436 20851 17440
rect 20787 17380 20791 17436
rect 20791 17380 20847 17436
rect 20847 17380 20851 17436
rect 20787 17376 20851 17380
rect 3401 16892 3465 16896
rect 3401 16836 3405 16892
rect 3405 16836 3461 16892
rect 3461 16836 3465 16892
rect 3401 16832 3465 16836
rect 3481 16892 3545 16896
rect 3481 16836 3485 16892
rect 3485 16836 3541 16892
rect 3541 16836 3545 16892
rect 3481 16832 3545 16836
rect 3561 16892 3625 16896
rect 3561 16836 3565 16892
rect 3565 16836 3621 16892
rect 3621 16836 3625 16892
rect 3561 16832 3625 16836
rect 3641 16892 3705 16896
rect 3641 16836 3645 16892
rect 3645 16836 3701 16892
rect 3701 16836 3705 16892
rect 3641 16832 3705 16836
rect 8300 16892 8364 16896
rect 8300 16836 8304 16892
rect 8304 16836 8360 16892
rect 8360 16836 8364 16892
rect 8300 16832 8364 16836
rect 8380 16892 8444 16896
rect 8380 16836 8384 16892
rect 8384 16836 8440 16892
rect 8440 16836 8444 16892
rect 8380 16832 8444 16836
rect 8460 16892 8524 16896
rect 8460 16836 8464 16892
rect 8464 16836 8520 16892
rect 8520 16836 8524 16892
rect 8460 16832 8524 16836
rect 8540 16892 8604 16896
rect 8540 16836 8544 16892
rect 8544 16836 8600 16892
rect 8600 16836 8604 16892
rect 8540 16832 8604 16836
rect 13199 16892 13263 16896
rect 13199 16836 13203 16892
rect 13203 16836 13259 16892
rect 13259 16836 13263 16892
rect 13199 16832 13263 16836
rect 13279 16892 13343 16896
rect 13279 16836 13283 16892
rect 13283 16836 13339 16892
rect 13339 16836 13343 16892
rect 13279 16832 13343 16836
rect 13359 16892 13423 16896
rect 13359 16836 13363 16892
rect 13363 16836 13419 16892
rect 13419 16836 13423 16892
rect 13359 16832 13423 16836
rect 13439 16892 13503 16896
rect 13439 16836 13443 16892
rect 13443 16836 13499 16892
rect 13499 16836 13503 16892
rect 13439 16832 13503 16836
rect 18098 16892 18162 16896
rect 18098 16836 18102 16892
rect 18102 16836 18158 16892
rect 18158 16836 18162 16892
rect 18098 16832 18162 16836
rect 18178 16892 18242 16896
rect 18178 16836 18182 16892
rect 18182 16836 18238 16892
rect 18238 16836 18242 16892
rect 18178 16832 18242 16836
rect 18258 16892 18322 16896
rect 18258 16836 18262 16892
rect 18262 16836 18318 16892
rect 18318 16836 18322 16892
rect 18258 16832 18322 16836
rect 18338 16892 18402 16896
rect 18338 16836 18342 16892
rect 18342 16836 18398 16892
rect 18398 16836 18402 16892
rect 18338 16832 18402 16836
rect 5850 16348 5914 16352
rect 5850 16292 5854 16348
rect 5854 16292 5910 16348
rect 5910 16292 5914 16348
rect 5850 16288 5914 16292
rect 5930 16348 5994 16352
rect 5930 16292 5934 16348
rect 5934 16292 5990 16348
rect 5990 16292 5994 16348
rect 5930 16288 5994 16292
rect 6010 16348 6074 16352
rect 6010 16292 6014 16348
rect 6014 16292 6070 16348
rect 6070 16292 6074 16348
rect 6010 16288 6074 16292
rect 6090 16348 6154 16352
rect 6090 16292 6094 16348
rect 6094 16292 6150 16348
rect 6150 16292 6154 16348
rect 6090 16288 6154 16292
rect 10749 16348 10813 16352
rect 10749 16292 10753 16348
rect 10753 16292 10809 16348
rect 10809 16292 10813 16348
rect 10749 16288 10813 16292
rect 10829 16348 10893 16352
rect 10829 16292 10833 16348
rect 10833 16292 10889 16348
rect 10889 16292 10893 16348
rect 10829 16288 10893 16292
rect 10909 16348 10973 16352
rect 10909 16292 10913 16348
rect 10913 16292 10969 16348
rect 10969 16292 10973 16348
rect 10909 16288 10973 16292
rect 10989 16348 11053 16352
rect 10989 16292 10993 16348
rect 10993 16292 11049 16348
rect 11049 16292 11053 16348
rect 10989 16288 11053 16292
rect 15648 16348 15712 16352
rect 15648 16292 15652 16348
rect 15652 16292 15708 16348
rect 15708 16292 15712 16348
rect 15648 16288 15712 16292
rect 15728 16348 15792 16352
rect 15728 16292 15732 16348
rect 15732 16292 15788 16348
rect 15788 16292 15792 16348
rect 15728 16288 15792 16292
rect 15808 16348 15872 16352
rect 15808 16292 15812 16348
rect 15812 16292 15868 16348
rect 15868 16292 15872 16348
rect 15808 16288 15872 16292
rect 15888 16348 15952 16352
rect 15888 16292 15892 16348
rect 15892 16292 15948 16348
rect 15948 16292 15952 16348
rect 15888 16288 15952 16292
rect 20547 16348 20611 16352
rect 20547 16292 20551 16348
rect 20551 16292 20607 16348
rect 20607 16292 20611 16348
rect 20547 16288 20611 16292
rect 20627 16348 20691 16352
rect 20627 16292 20631 16348
rect 20631 16292 20687 16348
rect 20687 16292 20691 16348
rect 20627 16288 20691 16292
rect 20707 16348 20771 16352
rect 20707 16292 20711 16348
rect 20711 16292 20767 16348
rect 20767 16292 20771 16348
rect 20707 16288 20771 16292
rect 20787 16348 20851 16352
rect 20787 16292 20791 16348
rect 20791 16292 20847 16348
rect 20847 16292 20851 16348
rect 20787 16288 20851 16292
rect 3401 15804 3465 15808
rect 3401 15748 3405 15804
rect 3405 15748 3461 15804
rect 3461 15748 3465 15804
rect 3401 15744 3465 15748
rect 3481 15804 3545 15808
rect 3481 15748 3485 15804
rect 3485 15748 3541 15804
rect 3541 15748 3545 15804
rect 3481 15744 3545 15748
rect 3561 15804 3625 15808
rect 3561 15748 3565 15804
rect 3565 15748 3621 15804
rect 3621 15748 3625 15804
rect 3561 15744 3625 15748
rect 3641 15804 3705 15808
rect 3641 15748 3645 15804
rect 3645 15748 3701 15804
rect 3701 15748 3705 15804
rect 3641 15744 3705 15748
rect 8300 15804 8364 15808
rect 8300 15748 8304 15804
rect 8304 15748 8360 15804
rect 8360 15748 8364 15804
rect 8300 15744 8364 15748
rect 8380 15804 8444 15808
rect 8380 15748 8384 15804
rect 8384 15748 8440 15804
rect 8440 15748 8444 15804
rect 8380 15744 8444 15748
rect 8460 15804 8524 15808
rect 8460 15748 8464 15804
rect 8464 15748 8520 15804
rect 8520 15748 8524 15804
rect 8460 15744 8524 15748
rect 8540 15804 8604 15808
rect 8540 15748 8544 15804
rect 8544 15748 8600 15804
rect 8600 15748 8604 15804
rect 8540 15744 8604 15748
rect 13199 15804 13263 15808
rect 13199 15748 13203 15804
rect 13203 15748 13259 15804
rect 13259 15748 13263 15804
rect 13199 15744 13263 15748
rect 13279 15804 13343 15808
rect 13279 15748 13283 15804
rect 13283 15748 13339 15804
rect 13339 15748 13343 15804
rect 13279 15744 13343 15748
rect 13359 15804 13423 15808
rect 13359 15748 13363 15804
rect 13363 15748 13419 15804
rect 13419 15748 13423 15804
rect 13359 15744 13423 15748
rect 13439 15804 13503 15808
rect 13439 15748 13443 15804
rect 13443 15748 13499 15804
rect 13499 15748 13503 15804
rect 13439 15744 13503 15748
rect 18098 15804 18162 15808
rect 18098 15748 18102 15804
rect 18102 15748 18158 15804
rect 18158 15748 18162 15804
rect 18098 15744 18162 15748
rect 18178 15804 18242 15808
rect 18178 15748 18182 15804
rect 18182 15748 18238 15804
rect 18238 15748 18242 15804
rect 18178 15744 18242 15748
rect 18258 15804 18322 15808
rect 18258 15748 18262 15804
rect 18262 15748 18318 15804
rect 18318 15748 18322 15804
rect 18258 15744 18322 15748
rect 18338 15804 18402 15808
rect 18338 15748 18342 15804
rect 18342 15748 18398 15804
rect 18398 15748 18402 15804
rect 18338 15744 18402 15748
rect 5850 15260 5914 15264
rect 5850 15204 5854 15260
rect 5854 15204 5910 15260
rect 5910 15204 5914 15260
rect 5850 15200 5914 15204
rect 5930 15260 5994 15264
rect 5930 15204 5934 15260
rect 5934 15204 5990 15260
rect 5990 15204 5994 15260
rect 5930 15200 5994 15204
rect 6010 15260 6074 15264
rect 6010 15204 6014 15260
rect 6014 15204 6070 15260
rect 6070 15204 6074 15260
rect 6010 15200 6074 15204
rect 6090 15260 6154 15264
rect 6090 15204 6094 15260
rect 6094 15204 6150 15260
rect 6150 15204 6154 15260
rect 6090 15200 6154 15204
rect 10749 15260 10813 15264
rect 10749 15204 10753 15260
rect 10753 15204 10809 15260
rect 10809 15204 10813 15260
rect 10749 15200 10813 15204
rect 10829 15260 10893 15264
rect 10829 15204 10833 15260
rect 10833 15204 10889 15260
rect 10889 15204 10893 15260
rect 10829 15200 10893 15204
rect 10909 15260 10973 15264
rect 10909 15204 10913 15260
rect 10913 15204 10969 15260
rect 10969 15204 10973 15260
rect 10909 15200 10973 15204
rect 10989 15260 11053 15264
rect 10989 15204 10993 15260
rect 10993 15204 11049 15260
rect 11049 15204 11053 15260
rect 10989 15200 11053 15204
rect 15648 15260 15712 15264
rect 15648 15204 15652 15260
rect 15652 15204 15708 15260
rect 15708 15204 15712 15260
rect 15648 15200 15712 15204
rect 15728 15260 15792 15264
rect 15728 15204 15732 15260
rect 15732 15204 15788 15260
rect 15788 15204 15792 15260
rect 15728 15200 15792 15204
rect 15808 15260 15872 15264
rect 15808 15204 15812 15260
rect 15812 15204 15868 15260
rect 15868 15204 15872 15260
rect 15808 15200 15872 15204
rect 15888 15260 15952 15264
rect 15888 15204 15892 15260
rect 15892 15204 15948 15260
rect 15948 15204 15952 15260
rect 15888 15200 15952 15204
rect 20547 15260 20611 15264
rect 20547 15204 20551 15260
rect 20551 15204 20607 15260
rect 20607 15204 20611 15260
rect 20547 15200 20611 15204
rect 20627 15260 20691 15264
rect 20627 15204 20631 15260
rect 20631 15204 20687 15260
rect 20687 15204 20691 15260
rect 20627 15200 20691 15204
rect 20707 15260 20771 15264
rect 20707 15204 20711 15260
rect 20711 15204 20767 15260
rect 20767 15204 20771 15260
rect 20707 15200 20771 15204
rect 20787 15260 20851 15264
rect 20787 15204 20791 15260
rect 20791 15204 20847 15260
rect 20847 15204 20851 15260
rect 20787 15200 20851 15204
rect 3401 14716 3465 14720
rect 3401 14660 3405 14716
rect 3405 14660 3461 14716
rect 3461 14660 3465 14716
rect 3401 14656 3465 14660
rect 3481 14716 3545 14720
rect 3481 14660 3485 14716
rect 3485 14660 3541 14716
rect 3541 14660 3545 14716
rect 3481 14656 3545 14660
rect 3561 14716 3625 14720
rect 3561 14660 3565 14716
rect 3565 14660 3621 14716
rect 3621 14660 3625 14716
rect 3561 14656 3625 14660
rect 3641 14716 3705 14720
rect 3641 14660 3645 14716
rect 3645 14660 3701 14716
rect 3701 14660 3705 14716
rect 3641 14656 3705 14660
rect 8300 14716 8364 14720
rect 8300 14660 8304 14716
rect 8304 14660 8360 14716
rect 8360 14660 8364 14716
rect 8300 14656 8364 14660
rect 8380 14716 8444 14720
rect 8380 14660 8384 14716
rect 8384 14660 8440 14716
rect 8440 14660 8444 14716
rect 8380 14656 8444 14660
rect 8460 14716 8524 14720
rect 8460 14660 8464 14716
rect 8464 14660 8520 14716
rect 8520 14660 8524 14716
rect 8460 14656 8524 14660
rect 8540 14716 8604 14720
rect 8540 14660 8544 14716
rect 8544 14660 8600 14716
rect 8600 14660 8604 14716
rect 8540 14656 8604 14660
rect 13199 14716 13263 14720
rect 13199 14660 13203 14716
rect 13203 14660 13259 14716
rect 13259 14660 13263 14716
rect 13199 14656 13263 14660
rect 13279 14716 13343 14720
rect 13279 14660 13283 14716
rect 13283 14660 13339 14716
rect 13339 14660 13343 14716
rect 13279 14656 13343 14660
rect 13359 14716 13423 14720
rect 13359 14660 13363 14716
rect 13363 14660 13419 14716
rect 13419 14660 13423 14716
rect 13359 14656 13423 14660
rect 13439 14716 13503 14720
rect 13439 14660 13443 14716
rect 13443 14660 13499 14716
rect 13499 14660 13503 14716
rect 13439 14656 13503 14660
rect 18098 14716 18162 14720
rect 18098 14660 18102 14716
rect 18102 14660 18158 14716
rect 18158 14660 18162 14716
rect 18098 14656 18162 14660
rect 18178 14716 18242 14720
rect 18178 14660 18182 14716
rect 18182 14660 18238 14716
rect 18238 14660 18242 14716
rect 18178 14656 18242 14660
rect 18258 14716 18322 14720
rect 18258 14660 18262 14716
rect 18262 14660 18318 14716
rect 18318 14660 18322 14716
rect 18258 14656 18322 14660
rect 18338 14716 18402 14720
rect 18338 14660 18342 14716
rect 18342 14660 18398 14716
rect 18398 14660 18402 14716
rect 18338 14656 18402 14660
rect 5850 14172 5914 14176
rect 5850 14116 5854 14172
rect 5854 14116 5910 14172
rect 5910 14116 5914 14172
rect 5850 14112 5914 14116
rect 5930 14172 5994 14176
rect 5930 14116 5934 14172
rect 5934 14116 5990 14172
rect 5990 14116 5994 14172
rect 5930 14112 5994 14116
rect 6010 14172 6074 14176
rect 6010 14116 6014 14172
rect 6014 14116 6070 14172
rect 6070 14116 6074 14172
rect 6010 14112 6074 14116
rect 6090 14172 6154 14176
rect 6090 14116 6094 14172
rect 6094 14116 6150 14172
rect 6150 14116 6154 14172
rect 6090 14112 6154 14116
rect 10749 14172 10813 14176
rect 10749 14116 10753 14172
rect 10753 14116 10809 14172
rect 10809 14116 10813 14172
rect 10749 14112 10813 14116
rect 10829 14172 10893 14176
rect 10829 14116 10833 14172
rect 10833 14116 10889 14172
rect 10889 14116 10893 14172
rect 10829 14112 10893 14116
rect 10909 14172 10973 14176
rect 10909 14116 10913 14172
rect 10913 14116 10969 14172
rect 10969 14116 10973 14172
rect 10909 14112 10973 14116
rect 10989 14172 11053 14176
rect 10989 14116 10993 14172
rect 10993 14116 11049 14172
rect 11049 14116 11053 14172
rect 10989 14112 11053 14116
rect 15648 14172 15712 14176
rect 15648 14116 15652 14172
rect 15652 14116 15708 14172
rect 15708 14116 15712 14172
rect 15648 14112 15712 14116
rect 15728 14172 15792 14176
rect 15728 14116 15732 14172
rect 15732 14116 15788 14172
rect 15788 14116 15792 14172
rect 15728 14112 15792 14116
rect 15808 14172 15872 14176
rect 15808 14116 15812 14172
rect 15812 14116 15868 14172
rect 15868 14116 15872 14172
rect 15808 14112 15872 14116
rect 15888 14172 15952 14176
rect 15888 14116 15892 14172
rect 15892 14116 15948 14172
rect 15948 14116 15952 14172
rect 15888 14112 15952 14116
rect 20547 14172 20611 14176
rect 20547 14116 20551 14172
rect 20551 14116 20607 14172
rect 20607 14116 20611 14172
rect 20547 14112 20611 14116
rect 20627 14172 20691 14176
rect 20627 14116 20631 14172
rect 20631 14116 20687 14172
rect 20687 14116 20691 14172
rect 20627 14112 20691 14116
rect 20707 14172 20771 14176
rect 20707 14116 20711 14172
rect 20711 14116 20767 14172
rect 20767 14116 20771 14172
rect 20707 14112 20771 14116
rect 20787 14172 20851 14176
rect 20787 14116 20791 14172
rect 20791 14116 20847 14172
rect 20847 14116 20851 14172
rect 20787 14112 20851 14116
rect 3401 13628 3465 13632
rect 3401 13572 3405 13628
rect 3405 13572 3461 13628
rect 3461 13572 3465 13628
rect 3401 13568 3465 13572
rect 3481 13628 3545 13632
rect 3481 13572 3485 13628
rect 3485 13572 3541 13628
rect 3541 13572 3545 13628
rect 3481 13568 3545 13572
rect 3561 13628 3625 13632
rect 3561 13572 3565 13628
rect 3565 13572 3621 13628
rect 3621 13572 3625 13628
rect 3561 13568 3625 13572
rect 3641 13628 3705 13632
rect 3641 13572 3645 13628
rect 3645 13572 3701 13628
rect 3701 13572 3705 13628
rect 3641 13568 3705 13572
rect 8300 13628 8364 13632
rect 8300 13572 8304 13628
rect 8304 13572 8360 13628
rect 8360 13572 8364 13628
rect 8300 13568 8364 13572
rect 8380 13628 8444 13632
rect 8380 13572 8384 13628
rect 8384 13572 8440 13628
rect 8440 13572 8444 13628
rect 8380 13568 8444 13572
rect 8460 13628 8524 13632
rect 8460 13572 8464 13628
rect 8464 13572 8520 13628
rect 8520 13572 8524 13628
rect 8460 13568 8524 13572
rect 8540 13628 8604 13632
rect 8540 13572 8544 13628
rect 8544 13572 8600 13628
rect 8600 13572 8604 13628
rect 8540 13568 8604 13572
rect 13199 13628 13263 13632
rect 13199 13572 13203 13628
rect 13203 13572 13259 13628
rect 13259 13572 13263 13628
rect 13199 13568 13263 13572
rect 13279 13628 13343 13632
rect 13279 13572 13283 13628
rect 13283 13572 13339 13628
rect 13339 13572 13343 13628
rect 13279 13568 13343 13572
rect 13359 13628 13423 13632
rect 13359 13572 13363 13628
rect 13363 13572 13419 13628
rect 13419 13572 13423 13628
rect 13359 13568 13423 13572
rect 13439 13628 13503 13632
rect 13439 13572 13443 13628
rect 13443 13572 13499 13628
rect 13499 13572 13503 13628
rect 13439 13568 13503 13572
rect 18098 13628 18162 13632
rect 18098 13572 18102 13628
rect 18102 13572 18158 13628
rect 18158 13572 18162 13628
rect 18098 13568 18162 13572
rect 18178 13628 18242 13632
rect 18178 13572 18182 13628
rect 18182 13572 18238 13628
rect 18238 13572 18242 13628
rect 18178 13568 18242 13572
rect 18258 13628 18322 13632
rect 18258 13572 18262 13628
rect 18262 13572 18318 13628
rect 18318 13572 18322 13628
rect 18258 13568 18322 13572
rect 18338 13628 18402 13632
rect 18338 13572 18342 13628
rect 18342 13572 18398 13628
rect 18398 13572 18402 13628
rect 18338 13568 18402 13572
rect 5850 13084 5914 13088
rect 5850 13028 5854 13084
rect 5854 13028 5910 13084
rect 5910 13028 5914 13084
rect 5850 13024 5914 13028
rect 5930 13084 5994 13088
rect 5930 13028 5934 13084
rect 5934 13028 5990 13084
rect 5990 13028 5994 13084
rect 5930 13024 5994 13028
rect 6010 13084 6074 13088
rect 6010 13028 6014 13084
rect 6014 13028 6070 13084
rect 6070 13028 6074 13084
rect 6010 13024 6074 13028
rect 6090 13084 6154 13088
rect 6090 13028 6094 13084
rect 6094 13028 6150 13084
rect 6150 13028 6154 13084
rect 6090 13024 6154 13028
rect 10749 13084 10813 13088
rect 10749 13028 10753 13084
rect 10753 13028 10809 13084
rect 10809 13028 10813 13084
rect 10749 13024 10813 13028
rect 10829 13084 10893 13088
rect 10829 13028 10833 13084
rect 10833 13028 10889 13084
rect 10889 13028 10893 13084
rect 10829 13024 10893 13028
rect 10909 13084 10973 13088
rect 10909 13028 10913 13084
rect 10913 13028 10969 13084
rect 10969 13028 10973 13084
rect 10909 13024 10973 13028
rect 10989 13084 11053 13088
rect 10989 13028 10993 13084
rect 10993 13028 11049 13084
rect 11049 13028 11053 13084
rect 10989 13024 11053 13028
rect 15648 13084 15712 13088
rect 15648 13028 15652 13084
rect 15652 13028 15708 13084
rect 15708 13028 15712 13084
rect 15648 13024 15712 13028
rect 15728 13084 15792 13088
rect 15728 13028 15732 13084
rect 15732 13028 15788 13084
rect 15788 13028 15792 13084
rect 15728 13024 15792 13028
rect 15808 13084 15872 13088
rect 15808 13028 15812 13084
rect 15812 13028 15868 13084
rect 15868 13028 15872 13084
rect 15808 13024 15872 13028
rect 15888 13084 15952 13088
rect 15888 13028 15892 13084
rect 15892 13028 15948 13084
rect 15948 13028 15952 13084
rect 15888 13024 15952 13028
rect 20547 13084 20611 13088
rect 20547 13028 20551 13084
rect 20551 13028 20607 13084
rect 20607 13028 20611 13084
rect 20547 13024 20611 13028
rect 20627 13084 20691 13088
rect 20627 13028 20631 13084
rect 20631 13028 20687 13084
rect 20687 13028 20691 13084
rect 20627 13024 20691 13028
rect 20707 13084 20771 13088
rect 20707 13028 20711 13084
rect 20711 13028 20767 13084
rect 20767 13028 20771 13084
rect 20707 13024 20771 13028
rect 20787 13084 20851 13088
rect 20787 13028 20791 13084
rect 20791 13028 20847 13084
rect 20847 13028 20851 13084
rect 20787 13024 20851 13028
rect 3401 12540 3465 12544
rect 3401 12484 3405 12540
rect 3405 12484 3461 12540
rect 3461 12484 3465 12540
rect 3401 12480 3465 12484
rect 3481 12540 3545 12544
rect 3481 12484 3485 12540
rect 3485 12484 3541 12540
rect 3541 12484 3545 12540
rect 3481 12480 3545 12484
rect 3561 12540 3625 12544
rect 3561 12484 3565 12540
rect 3565 12484 3621 12540
rect 3621 12484 3625 12540
rect 3561 12480 3625 12484
rect 3641 12540 3705 12544
rect 3641 12484 3645 12540
rect 3645 12484 3701 12540
rect 3701 12484 3705 12540
rect 3641 12480 3705 12484
rect 8300 12540 8364 12544
rect 8300 12484 8304 12540
rect 8304 12484 8360 12540
rect 8360 12484 8364 12540
rect 8300 12480 8364 12484
rect 8380 12540 8444 12544
rect 8380 12484 8384 12540
rect 8384 12484 8440 12540
rect 8440 12484 8444 12540
rect 8380 12480 8444 12484
rect 8460 12540 8524 12544
rect 8460 12484 8464 12540
rect 8464 12484 8520 12540
rect 8520 12484 8524 12540
rect 8460 12480 8524 12484
rect 8540 12540 8604 12544
rect 8540 12484 8544 12540
rect 8544 12484 8600 12540
rect 8600 12484 8604 12540
rect 8540 12480 8604 12484
rect 13199 12540 13263 12544
rect 13199 12484 13203 12540
rect 13203 12484 13259 12540
rect 13259 12484 13263 12540
rect 13199 12480 13263 12484
rect 13279 12540 13343 12544
rect 13279 12484 13283 12540
rect 13283 12484 13339 12540
rect 13339 12484 13343 12540
rect 13279 12480 13343 12484
rect 13359 12540 13423 12544
rect 13359 12484 13363 12540
rect 13363 12484 13419 12540
rect 13419 12484 13423 12540
rect 13359 12480 13423 12484
rect 13439 12540 13503 12544
rect 13439 12484 13443 12540
rect 13443 12484 13499 12540
rect 13499 12484 13503 12540
rect 13439 12480 13503 12484
rect 18098 12540 18162 12544
rect 18098 12484 18102 12540
rect 18102 12484 18158 12540
rect 18158 12484 18162 12540
rect 18098 12480 18162 12484
rect 18178 12540 18242 12544
rect 18178 12484 18182 12540
rect 18182 12484 18238 12540
rect 18238 12484 18242 12540
rect 18178 12480 18242 12484
rect 18258 12540 18322 12544
rect 18258 12484 18262 12540
rect 18262 12484 18318 12540
rect 18318 12484 18322 12540
rect 18258 12480 18322 12484
rect 18338 12540 18402 12544
rect 18338 12484 18342 12540
rect 18342 12484 18398 12540
rect 18398 12484 18402 12540
rect 18338 12480 18402 12484
rect 5850 11996 5914 12000
rect 5850 11940 5854 11996
rect 5854 11940 5910 11996
rect 5910 11940 5914 11996
rect 5850 11936 5914 11940
rect 5930 11996 5994 12000
rect 5930 11940 5934 11996
rect 5934 11940 5990 11996
rect 5990 11940 5994 11996
rect 5930 11936 5994 11940
rect 6010 11996 6074 12000
rect 6010 11940 6014 11996
rect 6014 11940 6070 11996
rect 6070 11940 6074 11996
rect 6010 11936 6074 11940
rect 6090 11996 6154 12000
rect 6090 11940 6094 11996
rect 6094 11940 6150 11996
rect 6150 11940 6154 11996
rect 6090 11936 6154 11940
rect 10749 11996 10813 12000
rect 10749 11940 10753 11996
rect 10753 11940 10809 11996
rect 10809 11940 10813 11996
rect 10749 11936 10813 11940
rect 10829 11996 10893 12000
rect 10829 11940 10833 11996
rect 10833 11940 10889 11996
rect 10889 11940 10893 11996
rect 10829 11936 10893 11940
rect 10909 11996 10973 12000
rect 10909 11940 10913 11996
rect 10913 11940 10969 11996
rect 10969 11940 10973 11996
rect 10909 11936 10973 11940
rect 10989 11996 11053 12000
rect 10989 11940 10993 11996
rect 10993 11940 11049 11996
rect 11049 11940 11053 11996
rect 10989 11936 11053 11940
rect 15648 11996 15712 12000
rect 15648 11940 15652 11996
rect 15652 11940 15708 11996
rect 15708 11940 15712 11996
rect 15648 11936 15712 11940
rect 15728 11996 15792 12000
rect 15728 11940 15732 11996
rect 15732 11940 15788 11996
rect 15788 11940 15792 11996
rect 15728 11936 15792 11940
rect 15808 11996 15872 12000
rect 15808 11940 15812 11996
rect 15812 11940 15868 11996
rect 15868 11940 15872 11996
rect 15808 11936 15872 11940
rect 15888 11996 15952 12000
rect 15888 11940 15892 11996
rect 15892 11940 15948 11996
rect 15948 11940 15952 11996
rect 15888 11936 15952 11940
rect 20547 11996 20611 12000
rect 20547 11940 20551 11996
rect 20551 11940 20607 11996
rect 20607 11940 20611 11996
rect 20547 11936 20611 11940
rect 20627 11996 20691 12000
rect 20627 11940 20631 11996
rect 20631 11940 20687 11996
rect 20687 11940 20691 11996
rect 20627 11936 20691 11940
rect 20707 11996 20771 12000
rect 20707 11940 20711 11996
rect 20711 11940 20767 11996
rect 20767 11940 20771 11996
rect 20707 11936 20771 11940
rect 20787 11996 20851 12000
rect 20787 11940 20791 11996
rect 20791 11940 20847 11996
rect 20847 11940 20851 11996
rect 20787 11936 20851 11940
rect 3401 11452 3465 11456
rect 3401 11396 3405 11452
rect 3405 11396 3461 11452
rect 3461 11396 3465 11452
rect 3401 11392 3465 11396
rect 3481 11452 3545 11456
rect 3481 11396 3485 11452
rect 3485 11396 3541 11452
rect 3541 11396 3545 11452
rect 3481 11392 3545 11396
rect 3561 11452 3625 11456
rect 3561 11396 3565 11452
rect 3565 11396 3621 11452
rect 3621 11396 3625 11452
rect 3561 11392 3625 11396
rect 3641 11452 3705 11456
rect 3641 11396 3645 11452
rect 3645 11396 3701 11452
rect 3701 11396 3705 11452
rect 3641 11392 3705 11396
rect 8300 11452 8364 11456
rect 8300 11396 8304 11452
rect 8304 11396 8360 11452
rect 8360 11396 8364 11452
rect 8300 11392 8364 11396
rect 8380 11452 8444 11456
rect 8380 11396 8384 11452
rect 8384 11396 8440 11452
rect 8440 11396 8444 11452
rect 8380 11392 8444 11396
rect 8460 11452 8524 11456
rect 8460 11396 8464 11452
rect 8464 11396 8520 11452
rect 8520 11396 8524 11452
rect 8460 11392 8524 11396
rect 8540 11452 8604 11456
rect 8540 11396 8544 11452
rect 8544 11396 8600 11452
rect 8600 11396 8604 11452
rect 8540 11392 8604 11396
rect 13199 11452 13263 11456
rect 13199 11396 13203 11452
rect 13203 11396 13259 11452
rect 13259 11396 13263 11452
rect 13199 11392 13263 11396
rect 13279 11452 13343 11456
rect 13279 11396 13283 11452
rect 13283 11396 13339 11452
rect 13339 11396 13343 11452
rect 13279 11392 13343 11396
rect 13359 11452 13423 11456
rect 13359 11396 13363 11452
rect 13363 11396 13419 11452
rect 13419 11396 13423 11452
rect 13359 11392 13423 11396
rect 13439 11452 13503 11456
rect 13439 11396 13443 11452
rect 13443 11396 13499 11452
rect 13499 11396 13503 11452
rect 13439 11392 13503 11396
rect 18098 11452 18162 11456
rect 18098 11396 18102 11452
rect 18102 11396 18158 11452
rect 18158 11396 18162 11452
rect 18098 11392 18162 11396
rect 18178 11452 18242 11456
rect 18178 11396 18182 11452
rect 18182 11396 18238 11452
rect 18238 11396 18242 11452
rect 18178 11392 18242 11396
rect 18258 11452 18322 11456
rect 18258 11396 18262 11452
rect 18262 11396 18318 11452
rect 18318 11396 18322 11452
rect 18258 11392 18322 11396
rect 18338 11452 18402 11456
rect 18338 11396 18342 11452
rect 18342 11396 18398 11452
rect 18398 11396 18402 11452
rect 18338 11392 18402 11396
rect 5850 10908 5914 10912
rect 5850 10852 5854 10908
rect 5854 10852 5910 10908
rect 5910 10852 5914 10908
rect 5850 10848 5914 10852
rect 5930 10908 5994 10912
rect 5930 10852 5934 10908
rect 5934 10852 5990 10908
rect 5990 10852 5994 10908
rect 5930 10848 5994 10852
rect 6010 10908 6074 10912
rect 6010 10852 6014 10908
rect 6014 10852 6070 10908
rect 6070 10852 6074 10908
rect 6010 10848 6074 10852
rect 6090 10908 6154 10912
rect 6090 10852 6094 10908
rect 6094 10852 6150 10908
rect 6150 10852 6154 10908
rect 6090 10848 6154 10852
rect 10749 10908 10813 10912
rect 10749 10852 10753 10908
rect 10753 10852 10809 10908
rect 10809 10852 10813 10908
rect 10749 10848 10813 10852
rect 10829 10908 10893 10912
rect 10829 10852 10833 10908
rect 10833 10852 10889 10908
rect 10889 10852 10893 10908
rect 10829 10848 10893 10852
rect 10909 10908 10973 10912
rect 10909 10852 10913 10908
rect 10913 10852 10969 10908
rect 10969 10852 10973 10908
rect 10909 10848 10973 10852
rect 10989 10908 11053 10912
rect 10989 10852 10993 10908
rect 10993 10852 11049 10908
rect 11049 10852 11053 10908
rect 10989 10848 11053 10852
rect 15648 10908 15712 10912
rect 15648 10852 15652 10908
rect 15652 10852 15708 10908
rect 15708 10852 15712 10908
rect 15648 10848 15712 10852
rect 15728 10908 15792 10912
rect 15728 10852 15732 10908
rect 15732 10852 15788 10908
rect 15788 10852 15792 10908
rect 15728 10848 15792 10852
rect 15808 10908 15872 10912
rect 15808 10852 15812 10908
rect 15812 10852 15868 10908
rect 15868 10852 15872 10908
rect 15808 10848 15872 10852
rect 15888 10908 15952 10912
rect 15888 10852 15892 10908
rect 15892 10852 15948 10908
rect 15948 10852 15952 10908
rect 15888 10848 15952 10852
rect 20547 10908 20611 10912
rect 20547 10852 20551 10908
rect 20551 10852 20607 10908
rect 20607 10852 20611 10908
rect 20547 10848 20611 10852
rect 20627 10908 20691 10912
rect 20627 10852 20631 10908
rect 20631 10852 20687 10908
rect 20687 10852 20691 10908
rect 20627 10848 20691 10852
rect 20707 10908 20771 10912
rect 20707 10852 20711 10908
rect 20711 10852 20767 10908
rect 20767 10852 20771 10908
rect 20707 10848 20771 10852
rect 20787 10908 20851 10912
rect 20787 10852 20791 10908
rect 20791 10852 20847 10908
rect 20847 10852 20851 10908
rect 20787 10848 20851 10852
rect 3401 10364 3465 10368
rect 3401 10308 3405 10364
rect 3405 10308 3461 10364
rect 3461 10308 3465 10364
rect 3401 10304 3465 10308
rect 3481 10364 3545 10368
rect 3481 10308 3485 10364
rect 3485 10308 3541 10364
rect 3541 10308 3545 10364
rect 3481 10304 3545 10308
rect 3561 10364 3625 10368
rect 3561 10308 3565 10364
rect 3565 10308 3621 10364
rect 3621 10308 3625 10364
rect 3561 10304 3625 10308
rect 3641 10364 3705 10368
rect 3641 10308 3645 10364
rect 3645 10308 3701 10364
rect 3701 10308 3705 10364
rect 3641 10304 3705 10308
rect 8300 10364 8364 10368
rect 8300 10308 8304 10364
rect 8304 10308 8360 10364
rect 8360 10308 8364 10364
rect 8300 10304 8364 10308
rect 8380 10364 8444 10368
rect 8380 10308 8384 10364
rect 8384 10308 8440 10364
rect 8440 10308 8444 10364
rect 8380 10304 8444 10308
rect 8460 10364 8524 10368
rect 8460 10308 8464 10364
rect 8464 10308 8520 10364
rect 8520 10308 8524 10364
rect 8460 10304 8524 10308
rect 8540 10364 8604 10368
rect 8540 10308 8544 10364
rect 8544 10308 8600 10364
rect 8600 10308 8604 10364
rect 8540 10304 8604 10308
rect 13199 10364 13263 10368
rect 13199 10308 13203 10364
rect 13203 10308 13259 10364
rect 13259 10308 13263 10364
rect 13199 10304 13263 10308
rect 13279 10364 13343 10368
rect 13279 10308 13283 10364
rect 13283 10308 13339 10364
rect 13339 10308 13343 10364
rect 13279 10304 13343 10308
rect 13359 10364 13423 10368
rect 13359 10308 13363 10364
rect 13363 10308 13419 10364
rect 13419 10308 13423 10364
rect 13359 10304 13423 10308
rect 13439 10364 13503 10368
rect 13439 10308 13443 10364
rect 13443 10308 13499 10364
rect 13499 10308 13503 10364
rect 13439 10304 13503 10308
rect 18098 10364 18162 10368
rect 18098 10308 18102 10364
rect 18102 10308 18158 10364
rect 18158 10308 18162 10364
rect 18098 10304 18162 10308
rect 18178 10364 18242 10368
rect 18178 10308 18182 10364
rect 18182 10308 18238 10364
rect 18238 10308 18242 10364
rect 18178 10304 18242 10308
rect 18258 10364 18322 10368
rect 18258 10308 18262 10364
rect 18262 10308 18318 10364
rect 18318 10308 18322 10364
rect 18258 10304 18322 10308
rect 18338 10364 18402 10368
rect 18338 10308 18342 10364
rect 18342 10308 18398 10364
rect 18398 10308 18402 10364
rect 18338 10304 18402 10308
rect 5850 9820 5914 9824
rect 5850 9764 5854 9820
rect 5854 9764 5910 9820
rect 5910 9764 5914 9820
rect 5850 9760 5914 9764
rect 5930 9820 5994 9824
rect 5930 9764 5934 9820
rect 5934 9764 5990 9820
rect 5990 9764 5994 9820
rect 5930 9760 5994 9764
rect 6010 9820 6074 9824
rect 6010 9764 6014 9820
rect 6014 9764 6070 9820
rect 6070 9764 6074 9820
rect 6010 9760 6074 9764
rect 6090 9820 6154 9824
rect 6090 9764 6094 9820
rect 6094 9764 6150 9820
rect 6150 9764 6154 9820
rect 6090 9760 6154 9764
rect 10749 9820 10813 9824
rect 10749 9764 10753 9820
rect 10753 9764 10809 9820
rect 10809 9764 10813 9820
rect 10749 9760 10813 9764
rect 10829 9820 10893 9824
rect 10829 9764 10833 9820
rect 10833 9764 10889 9820
rect 10889 9764 10893 9820
rect 10829 9760 10893 9764
rect 10909 9820 10973 9824
rect 10909 9764 10913 9820
rect 10913 9764 10969 9820
rect 10969 9764 10973 9820
rect 10909 9760 10973 9764
rect 10989 9820 11053 9824
rect 10989 9764 10993 9820
rect 10993 9764 11049 9820
rect 11049 9764 11053 9820
rect 10989 9760 11053 9764
rect 15648 9820 15712 9824
rect 15648 9764 15652 9820
rect 15652 9764 15708 9820
rect 15708 9764 15712 9820
rect 15648 9760 15712 9764
rect 15728 9820 15792 9824
rect 15728 9764 15732 9820
rect 15732 9764 15788 9820
rect 15788 9764 15792 9820
rect 15728 9760 15792 9764
rect 15808 9820 15872 9824
rect 15808 9764 15812 9820
rect 15812 9764 15868 9820
rect 15868 9764 15872 9820
rect 15808 9760 15872 9764
rect 15888 9820 15952 9824
rect 15888 9764 15892 9820
rect 15892 9764 15948 9820
rect 15948 9764 15952 9820
rect 15888 9760 15952 9764
rect 20547 9820 20611 9824
rect 20547 9764 20551 9820
rect 20551 9764 20607 9820
rect 20607 9764 20611 9820
rect 20547 9760 20611 9764
rect 20627 9820 20691 9824
rect 20627 9764 20631 9820
rect 20631 9764 20687 9820
rect 20687 9764 20691 9820
rect 20627 9760 20691 9764
rect 20707 9820 20771 9824
rect 20707 9764 20711 9820
rect 20711 9764 20767 9820
rect 20767 9764 20771 9820
rect 20707 9760 20771 9764
rect 20787 9820 20851 9824
rect 20787 9764 20791 9820
rect 20791 9764 20847 9820
rect 20847 9764 20851 9820
rect 20787 9760 20851 9764
rect 3401 9276 3465 9280
rect 3401 9220 3405 9276
rect 3405 9220 3461 9276
rect 3461 9220 3465 9276
rect 3401 9216 3465 9220
rect 3481 9276 3545 9280
rect 3481 9220 3485 9276
rect 3485 9220 3541 9276
rect 3541 9220 3545 9276
rect 3481 9216 3545 9220
rect 3561 9276 3625 9280
rect 3561 9220 3565 9276
rect 3565 9220 3621 9276
rect 3621 9220 3625 9276
rect 3561 9216 3625 9220
rect 3641 9276 3705 9280
rect 3641 9220 3645 9276
rect 3645 9220 3701 9276
rect 3701 9220 3705 9276
rect 3641 9216 3705 9220
rect 8300 9276 8364 9280
rect 8300 9220 8304 9276
rect 8304 9220 8360 9276
rect 8360 9220 8364 9276
rect 8300 9216 8364 9220
rect 8380 9276 8444 9280
rect 8380 9220 8384 9276
rect 8384 9220 8440 9276
rect 8440 9220 8444 9276
rect 8380 9216 8444 9220
rect 8460 9276 8524 9280
rect 8460 9220 8464 9276
rect 8464 9220 8520 9276
rect 8520 9220 8524 9276
rect 8460 9216 8524 9220
rect 8540 9276 8604 9280
rect 8540 9220 8544 9276
rect 8544 9220 8600 9276
rect 8600 9220 8604 9276
rect 8540 9216 8604 9220
rect 13199 9276 13263 9280
rect 13199 9220 13203 9276
rect 13203 9220 13259 9276
rect 13259 9220 13263 9276
rect 13199 9216 13263 9220
rect 13279 9276 13343 9280
rect 13279 9220 13283 9276
rect 13283 9220 13339 9276
rect 13339 9220 13343 9276
rect 13279 9216 13343 9220
rect 13359 9276 13423 9280
rect 13359 9220 13363 9276
rect 13363 9220 13419 9276
rect 13419 9220 13423 9276
rect 13359 9216 13423 9220
rect 13439 9276 13503 9280
rect 13439 9220 13443 9276
rect 13443 9220 13499 9276
rect 13499 9220 13503 9276
rect 13439 9216 13503 9220
rect 18098 9276 18162 9280
rect 18098 9220 18102 9276
rect 18102 9220 18158 9276
rect 18158 9220 18162 9276
rect 18098 9216 18162 9220
rect 18178 9276 18242 9280
rect 18178 9220 18182 9276
rect 18182 9220 18238 9276
rect 18238 9220 18242 9276
rect 18178 9216 18242 9220
rect 18258 9276 18322 9280
rect 18258 9220 18262 9276
rect 18262 9220 18318 9276
rect 18318 9220 18322 9276
rect 18258 9216 18322 9220
rect 18338 9276 18402 9280
rect 18338 9220 18342 9276
rect 18342 9220 18398 9276
rect 18398 9220 18402 9276
rect 18338 9216 18402 9220
rect 5850 8732 5914 8736
rect 5850 8676 5854 8732
rect 5854 8676 5910 8732
rect 5910 8676 5914 8732
rect 5850 8672 5914 8676
rect 5930 8732 5994 8736
rect 5930 8676 5934 8732
rect 5934 8676 5990 8732
rect 5990 8676 5994 8732
rect 5930 8672 5994 8676
rect 6010 8732 6074 8736
rect 6010 8676 6014 8732
rect 6014 8676 6070 8732
rect 6070 8676 6074 8732
rect 6010 8672 6074 8676
rect 6090 8732 6154 8736
rect 6090 8676 6094 8732
rect 6094 8676 6150 8732
rect 6150 8676 6154 8732
rect 6090 8672 6154 8676
rect 10749 8732 10813 8736
rect 10749 8676 10753 8732
rect 10753 8676 10809 8732
rect 10809 8676 10813 8732
rect 10749 8672 10813 8676
rect 10829 8732 10893 8736
rect 10829 8676 10833 8732
rect 10833 8676 10889 8732
rect 10889 8676 10893 8732
rect 10829 8672 10893 8676
rect 10909 8732 10973 8736
rect 10909 8676 10913 8732
rect 10913 8676 10969 8732
rect 10969 8676 10973 8732
rect 10909 8672 10973 8676
rect 10989 8732 11053 8736
rect 10989 8676 10993 8732
rect 10993 8676 11049 8732
rect 11049 8676 11053 8732
rect 10989 8672 11053 8676
rect 15648 8732 15712 8736
rect 15648 8676 15652 8732
rect 15652 8676 15708 8732
rect 15708 8676 15712 8732
rect 15648 8672 15712 8676
rect 15728 8732 15792 8736
rect 15728 8676 15732 8732
rect 15732 8676 15788 8732
rect 15788 8676 15792 8732
rect 15728 8672 15792 8676
rect 15808 8732 15872 8736
rect 15808 8676 15812 8732
rect 15812 8676 15868 8732
rect 15868 8676 15872 8732
rect 15808 8672 15872 8676
rect 15888 8732 15952 8736
rect 15888 8676 15892 8732
rect 15892 8676 15948 8732
rect 15948 8676 15952 8732
rect 15888 8672 15952 8676
rect 20547 8732 20611 8736
rect 20547 8676 20551 8732
rect 20551 8676 20607 8732
rect 20607 8676 20611 8732
rect 20547 8672 20611 8676
rect 20627 8732 20691 8736
rect 20627 8676 20631 8732
rect 20631 8676 20687 8732
rect 20687 8676 20691 8732
rect 20627 8672 20691 8676
rect 20707 8732 20771 8736
rect 20707 8676 20711 8732
rect 20711 8676 20767 8732
rect 20767 8676 20771 8732
rect 20707 8672 20771 8676
rect 20787 8732 20851 8736
rect 20787 8676 20791 8732
rect 20791 8676 20847 8732
rect 20847 8676 20851 8732
rect 20787 8672 20851 8676
rect 3401 8188 3465 8192
rect 3401 8132 3405 8188
rect 3405 8132 3461 8188
rect 3461 8132 3465 8188
rect 3401 8128 3465 8132
rect 3481 8188 3545 8192
rect 3481 8132 3485 8188
rect 3485 8132 3541 8188
rect 3541 8132 3545 8188
rect 3481 8128 3545 8132
rect 3561 8188 3625 8192
rect 3561 8132 3565 8188
rect 3565 8132 3621 8188
rect 3621 8132 3625 8188
rect 3561 8128 3625 8132
rect 3641 8188 3705 8192
rect 3641 8132 3645 8188
rect 3645 8132 3701 8188
rect 3701 8132 3705 8188
rect 3641 8128 3705 8132
rect 8300 8188 8364 8192
rect 8300 8132 8304 8188
rect 8304 8132 8360 8188
rect 8360 8132 8364 8188
rect 8300 8128 8364 8132
rect 8380 8188 8444 8192
rect 8380 8132 8384 8188
rect 8384 8132 8440 8188
rect 8440 8132 8444 8188
rect 8380 8128 8444 8132
rect 8460 8188 8524 8192
rect 8460 8132 8464 8188
rect 8464 8132 8520 8188
rect 8520 8132 8524 8188
rect 8460 8128 8524 8132
rect 8540 8188 8604 8192
rect 8540 8132 8544 8188
rect 8544 8132 8600 8188
rect 8600 8132 8604 8188
rect 8540 8128 8604 8132
rect 13199 8188 13263 8192
rect 13199 8132 13203 8188
rect 13203 8132 13259 8188
rect 13259 8132 13263 8188
rect 13199 8128 13263 8132
rect 13279 8188 13343 8192
rect 13279 8132 13283 8188
rect 13283 8132 13339 8188
rect 13339 8132 13343 8188
rect 13279 8128 13343 8132
rect 13359 8188 13423 8192
rect 13359 8132 13363 8188
rect 13363 8132 13419 8188
rect 13419 8132 13423 8188
rect 13359 8128 13423 8132
rect 13439 8188 13503 8192
rect 13439 8132 13443 8188
rect 13443 8132 13499 8188
rect 13499 8132 13503 8188
rect 13439 8128 13503 8132
rect 18098 8188 18162 8192
rect 18098 8132 18102 8188
rect 18102 8132 18158 8188
rect 18158 8132 18162 8188
rect 18098 8128 18162 8132
rect 18178 8188 18242 8192
rect 18178 8132 18182 8188
rect 18182 8132 18238 8188
rect 18238 8132 18242 8188
rect 18178 8128 18242 8132
rect 18258 8188 18322 8192
rect 18258 8132 18262 8188
rect 18262 8132 18318 8188
rect 18318 8132 18322 8188
rect 18258 8128 18322 8132
rect 18338 8188 18402 8192
rect 18338 8132 18342 8188
rect 18342 8132 18398 8188
rect 18398 8132 18402 8188
rect 18338 8128 18402 8132
rect 5850 7644 5914 7648
rect 5850 7588 5854 7644
rect 5854 7588 5910 7644
rect 5910 7588 5914 7644
rect 5850 7584 5914 7588
rect 5930 7644 5994 7648
rect 5930 7588 5934 7644
rect 5934 7588 5990 7644
rect 5990 7588 5994 7644
rect 5930 7584 5994 7588
rect 6010 7644 6074 7648
rect 6010 7588 6014 7644
rect 6014 7588 6070 7644
rect 6070 7588 6074 7644
rect 6010 7584 6074 7588
rect 6090 7644 6154 7648
rect 6090 7588 6094 7644
rect 6094 7588 6150 7644
rect 6150 7588 6154 7644
rect 6090 7584 6154 7588
rect 10749 7644 10813 7648
rect 10749 7588 10753 7644
rect 10753 7588 10809 7644
rect 10809 7588 10813 7644
rect 10749 7584 10813 7588
rect 10829 7644 10893 7648
rect 10829 7588 10833 7644
rect 10833 7588 10889 7644
rect 10889 7588 10893 7644
rect 10829 7584 10893 7588
rect 10909 7644 10973 7648
rect 10909 7588 10913 7644
rect 10913 7588 10969 7644
rect 10969 7588 10973 7644
rect 10909 7584 10973 7588
rect 10989 7644 11053 7648
rect 10989 7588 10993 7644
rect 10993 7588 11049 7644
rect 11049 7588 11053 7644
rect 10989 7584 11053 7588
rect 15648 7644 15712 7648
rect 15648 7588 15652 7644
rect 15652 7588 15708 7644
rect 15708 7588 15712 7644
rect 15648 7584 15712 7588
rect 15728 7644 15792 7648
rect 15728 7588 15732 7644
rect 15732 7588 15788 7644
rect 15788 7588 15792 7644
rect 15728 7584 15792 7588
rect 15808 7644 15872 7648
rect 15808 7588 15812 7644
rect 15812 7588 15868 7644
rect 15868 7588 15872 7644
rect 15808 7584 15872 7588
rect 15888 7644 15952 7648
rect 15888 7588 15892 7644
rect 15892 7588 15948 7644
rect 15948 7588 15952 7644
rect 15888 7584 15952 7588
rect 20547 7644 20611 7648
rect 20547 7588 20551 7644
rect 20551 7588 20607 7644
rect 20607 7588 20611 7644
rect 20547 7584 20611 7588
rect 20627 7644 20691 7648
rect 20627 7588 20631 7644
rect 20631 7588 20687 7644
rect 20687 7588 20691 7644
rect 20627 7584 20691 7588
rect 20707 7644 20771 7648
rect 20707 7588 20711 7644
rect 20711 7588 20767 7644
rect 20767 7588 20771 7644
rect 20707 7584 20771 7588
rect 20787 7644 20851 7648
rect 20787 7588 20791 7644
rect 20791 7588 20847 7644
rect 20847 7588 20851 7644
rect 20787 7584 20851 7588
rect 3401 7100 3465 7104
rect 3401 7044 3405 7100
rect 3405 7044 3461 7100
rect 3461 7044 3465 7100
rect 3401 7040 3465 7044
rect 3481 7100 3545 7104
rect 3481 7044 3485 7100
rect 3485 7044 3541 7100
rect 3541 7044 3545 7100
rect 3481 7040 3545 7044
rect 3561 7100 3625 7104
rect 3561 7044 3565 7100
rect 3565 7044 3621 7100
rect 3621 7044 3625 7100
rect 3561 7040 3625 7044
rect 3641 7100 3705 7104
rect 3641 7044 3645 7100
rect 3645 7044 3701 7100
rect 3701 7044 3705 7100
rect 3641 7040 3705 7044
rect 8300 7100 8364 7104
rect 8300 7044 8304 7100
rect 8304 7044 8360 7100
rect 8360 7044 8364 7100
rect 8300 7040 8364 7044
rect 8380 7100 8444 7104
rect 8380 7044 8384 7100
rect 8384 7044 8440 7100
rect 8440 7044 8444 7100
rect 8380 7040 8444 7044
rect 8460 7100 8524 7104
rect 8460 7044 8464 7100
rect 8464 7044 8520 7100
rect 8520 7044 8524 7100
rect 8460 7040 8524 7044
rect 8540 7100 8604 7104
rect 8540 7044 8544 7100
rect 8544 7044 8600 7100
rect 8600 7044 8604 7100
rect 8540 7040 8604 7044
rect 13199 7100 13263 7104
rect 13199 7044 13203 7100
rect 13203 7044 13259 7100
rect 13259 7044 13263 7100
rect 13199 7040 13263 7044
rect 13279 7100 13343 7104
rect 13279 7044 13283 7100
rect 13283 7044 13339 7100
rect 13339 7044 13343 7100
rect 13279 7040 13343 7044
rect 13359 7100 13423 7104
rect 13359 7044 13363 7100
rect 13363 7044 13419 7100
rect 13419 7044 13423 7100
rect 13359 7040 13423 7044
rect 13439 7100 13503 7104
rect 13439 7044 13443 7100
rect 13443 7044 13499 7100
rect 13499 7044 13503 7100
rect 13439 7040 13503 7044
rect 18098 7100 18162 7104
rect 18098 7044 18102 7100
rect 18102 7044 18158 7100
rect 18158 7044 18162 7100
rect 18098 7040 18162 7044
rect 18178 7100 18242 7104
rect 18178 7044 18182 7100
rect 18182 7044 18238 7100
rect 18238 7044 18242 7100
rect 18178 7040 18242 7044
rect 18258 7100 18322 7104
rect 18258 7044 18262 7100
rect 18262 7044 18318 7100
rect 18318 7044 18322 7100
rect 18258 7040 18322 7044
rect 18338 7100 18402 7104
rect 18338 7044 18342 7100
rect 18342 7044 18398 7100
rect 18398 7044 18402 7100
rect 18338 7040 18402 7044
rect 5850 6556 5914 6560
rect 5850 6500 5854 6556
rect 5854 6500 5910 6556
rect 5910 6500 5914 6556
rect 5850 6496 5914 6500
rect 5930 6556 5994 6560
rect 5930 6500 5934 6556
rect 5934 6500 5990 6556
rect 5990 6500 5994 6556
rect 5930 6496 5994 6500
rect 6010 6556 6074 6560
rect 6010 6500 6014 6556
rect 6014 6500 6070 6556
rect 6070 6500 6074 6556
rect 6010 6496 6074 6500
rect 6090 6556 6154 6560
rect 6090 6500 6094 6556
rect 6094 6500 6150 6556
rect 6150 6500 6154 6556
rect 6090 6496 6154 6500
rect 10749 6556 10813 6560
rect 10749 6500 10753 6556
rect 10753 6500 10809 6556
rect 10809 6500 10813 6556
rect 10749 6496 10813 6500
rect 10829 6556 10893 6560
rect 10829 6500 10833 6556
rect 10833 6500 10889 6556
rect 10889 6500 10893 6556
rect 10829 6496 10893 6500
rect 10909 6556 10973 6560
rect 10909 6500 10913 6556
rect 10913 6500 10969 6556
rect 10969 6500 10973 6556
rect 10909 6496 10973 6500
rect 10989 6556 11053 6560
rect 10989 6500 10993 6556
rect 10993 6500 11049 6556
rect 11049 6500 11053 6556
rect 10989 6496 11053 6500
rect 15648 6556 15712 6560
rect 15648 6500 15652 6556
rect 15652 6500 15708 6556
rect 15708 6500 15712 6556
rect 15648 6496 15712 6500
rect 15728 6556 15792 6560
rect 15728 6500 15732 6556
rect 15732 6500 15788 6556
rect 15788 6500 15792 6556
rect 15728 6496 15792 6500
rect 15808 6556 15872 6560
rect 15808 6500 15812 6556
rect 15812 6500 15868 6556
rect 15868 6500 15872 6556
rect 15808 6496 15872 6500
rect 15888 6556 15952 6560
rect 15888 6500 15892 6556
rect 15892 6500 15948 6556
rect 15948 6500 15952 6556
rect 15888 6496 15952 6500
rect 20547 6556 20611 6560
rect 20547 6500 20551 6556
rect 20551 6500 20607 6556
rect 20607 6500 20611 6556
rect 20547 6496 20611 6500
rect 20627 6556 20691 6560
rect 20627 6500 20631 6556
rect 20631 6500 20687 6556
rect 20687 6500 20691 6556
rect 20627 6496 20691 6500
rect 20707 6556 20771 6560
rect 20707 6500 20711 6556
rect 20711 6500 20767 6556
rect 20767 6500 20771 6556
rect 20707 6496 20771 6500
rect 20787 6556 20851 6560
rect 20787 6500 20791 6556
rect 20791 6500 20847 6556
rect 20847 6500 20851 6556
rect 20787 6496 20851 6500
rect 3401 6012 3465 6016
rect 3401 5956 3405 6012
rect 3405 5956 3461 6012
rect 3461 5956 3465 6012
rect 3401 5952 3465 5956
rect 3481 6012 3545 6016
rect 3481 5956 3485 6012
rect 3485 5956 3541 6012
rect 3541 5956 3545 6012
rect 3481 5952 3545 5956
rect 3561 6012 3625 6016
rect 3561 5956 3565 6012
rect 3565 5956 3621 6012
rect 3621 5956 3625 6012
rect 3561 5952 3625 5956
rect 3641 6012 3705 6016
rect 3641 5956 3645 6012
rect 3645 5956 3701 6012
rect 3701 5956 3705 6012
rect 3641 5952 3705 5956
rect 8300 6012 8364 6016
rect 8300 5956 8304 6012
rect 8304 5956 8360 6012
rect 8360 5956 8364 6012
rect 8300 5952 8364 5956
rect 8380 6012 8444 6016
rect 8380 5956 8384 6012
rect 8384 5956 8440 6012
rect 8440 5956 8444 6012
rect 8380 5952 8444 5956
rect 8460 6012 8524 6016
rect 8460 5956 8464 6012
rect 8464 5956 8520 6012
rect 8520 5956 8524 6012
rect 8460 5952 8524 5956
rect 8540 6012 8604 6016
rect 8540 5956 8544 6012
rect 8544 5956 8600 6012
rect 8600 5956 8604 6012
rect 8540 5952 8604 5956
rect 13199 6012 13263 6016
rect 13199 5956 13203 6012
rect 13203 5956 13259 6012
rect 13259 5956 13263 6012
rect 13199 5952 13263 5956
rect 13279 6012 13343 6016
rect 13279 5956 13283 6012
rect 13283 5956 13339 6012
rect 13339 5956 13343 6012
rect 13279 5952 13343 5956
rect 13359 6012 13423 6016
rect 13359 5956 13363 6012
rect 13363 5956 13419 6012
rect 13419 5956 13423 6012
rect 13359 5952 13423 5956
rect 13439 6012 13503 6016
rect 13439 5956 13443 6012
rect 13443 5956 13499 6012
rect 13499 5956 13503 6012
rect 13439 5952 13503 5956
rect 18098 6012 18162 6016
rect 18098 5956 18102 6012
rect 18102 5956 18158 6012
rect 18158 5956 18162 6012
rect 18098 5952 18162 5956
rect 18178 6012 18242 6016
rect 18178 5956 18182 6012
rect 18182 5956 18238 6012
rect 18238 5956 18242 6012
rect 18178 5952 18242 5956
rect 18258 6012 18322 6016
rect 18258 5956 18262 6012
rect 18262 5956 18318 6012
rect 18318 5956 18322 6012
rect 18258 5952 18322 5956
rect 18338 6012 18402 6016
rect 18338 5956 18342 6012
rect 18342 5956 18398 6012
rect 18398 5956 18402 6012
rect 18338 5952 18402 5956
rect 5850 5468 5914 5472
rect 5850 5412 5854 5468
rect 5854 5412 5910 5468
rect 5910 5412 5914 5468
rect 5850 5408 5914 5412
rect 5930 5468 5994 5472
rect 5930 5412 5934 5468
rect 5934 5412 5990 5468
rect 5990 5412 5994 5468
rect 5930 5408 5994 5412
rect 6010 5468 6074 5472
rect 6010 5412 6014 5468
rect 6014 5412 6070 5468
rect 6070 5412 6074 5468
rect 6010 5408 6074 5412
rect 6090 5468 6154 5472
rect 6090 5412 6094 5468
rect 6094 5412 6150 5468
rect 6150 5412 6154 5468
rect 6090 5408 6154 5412
rect 10749 5468 10813 5472
rect 10749 5412 10753 5468
rect 10753 5412 10809 5468
rect 10809 5412 10813 5468
rect 10749 5408 10813 5412
rect 10829 5468 10893 5472
rect 10829 5412 10833 5468
rect 10833 5412 10889 5468
rect 10889 5412 10893 5468
rect 10829 5408 10893 5412
rect 10909 5468 10973 5472
rect 10909 5412 10913 5468
rect 10913 5412 10969 5468
rect 10969 5412 10973 5468
rect 10909 5408 10973 5412
rect 10989 5468 11053 5472
rect 10989 5412 10993 5468
rect 10993 5412 11049 5468
rect 11049 5412 11053 5468
rect 10989 5408 11053 5412
rect 15648 5468 15712 5472
rect 15648 5412 15652 5468
rect 15652 5412 15708 5468
rect 15708 5412 15712 5468
rect 15648 5408 15712 5412
rect 15728 5468 15792 5472
rect 15728 5412 15732 5468
rect 15732 5412 15788 5468
rect 15788 5412 15792 5468
rect 15728 5408 15792 5412
rect 15808 5468 15872 5472
rect 15808 5412 15812 5468
rect 15812 5412 15868 5468
rect 15868 5412 15872 5468
rect 15808 5408 15872 5412
rect 15888 5468 15952 5472
rect 15888 5412 15892 5468
rect 15892 5412 15948 5468
rect 15948 5412 15952 5468
rect 15888 5408 15952 5412
rect 20547 5468 20611 5472
rect 20547 5412 20551 5468
rect 20551 5412 20607 5468
rect 20607 5412 20611 5468
rect 20547 5408 20611 5412
rect 20627 5468 20691 5472
rect 20627 5412 20631 5468
rect 20631 5412 20687 5468
rect 20687 5412 20691 5468
rect 20627 5408 20691 5412
rect 20707 5468 20771 5472
rect 20707 5412 20711 5468
rect 20711 5412 20767 5468
rect 20767 5412 20771 5468
rect 20707 5408 20771 5412
rect 20787 5468 20851 5472
rect 20787 5412 20791 5468
rect 20791 5412 20847 5468
rect 20847 5412 20851 5468
rect 20787 5408 20851 5412
rect 3401 4924 3465 4928
rect 3401 4868 3405 4924
rect 3405 4868 3461 4924
rect 3461 4868 3465 4924
rect 3401 4864 3465 4868
rect 3481 4924 3545 4928
rect 3481 4868 3485 4924
rect 3485 4868 3541 4924
rect 3541 4868 3545 4924
rect 3481 4864 3545 4868
rect 3561 4924 3625 4928
rect 3561 4868 3565 4924
rect 3565 4868 3621 4924
rect 3621 4868 3625 4924
rect 3561 4864 3625 4868
rect 3641 4924 3705 4928
rect 3641 4868 3645 4924
rect 3645 4868 3701 4924
rect 3701 4868 3705 4924
rect 3641 4864 3705 4868
rect 8300 4924 8364 4928
rect 8300 4868 8304 4924
rect 8304 4868 8360 4924
rect 8360 4868 8364 4924
rect 8300 4864 8364 4868
rect 8380 4924 8444 4928
rect 8380 4868 8384 4924
rect 8384 4868 8440 4924
rect 8440 4868 8444 4924
rect 8380 4864 8444 4868
rect 8460 4924 8524 4928
rect 8460 4868 8464 4924
rect 8464 4868 8520 4924
rect 8520 4868 8524 4924
rect 8460 4864 8524 4868
rect 8540 4924 8604 4928
rect 8540 4868 8544 4924
rect 8544 4868 8600 4924
rect 8600 4868 8604 4924
rect 8540 4864 8604 4868
rect 13199 4924 13263 4928
rect 13199 4868 13203 4924
rect 13203 4868 13259 4924
rect 13259 4868 13263 4924
rect 13199 4864 13263 4868
rect 13279 4924 13343 4928
rect 13279 4868 13283 4924
rect 13283 4868 13339 4924
rect 13339 4868 13343 4924
rect 13279 4864 13343 4868
rect 13359 4924 13423 4928
rect 13359 4868 13363 4924
rect 13363 4868 13419 4924
rect 13419 4868 13423 4924
rect 13359 4864 13423 4868
rect 13439 4924 13503 4928
rect 13439 4868 13443 4924
rect 13443 4868 13499 4924
rect 13499 4868 13503 4924
rect 13439 4864 13503 4868
rect 18098 4924 18162 4928
rect 18098 4868 18102 4924
rect 18102 4868 18158 4924
rect 18158 4868 18162 4924
rect 18098 4864 18162 4868
rect 18178 4924 18242 4928
rect 18178 4868 18182 4924
rect 18182 4868 18238 4924
rect 18238 4868 18242 4924
rect 18178 4864 18242 4868
rect 18258 4924 18322 4928
rect 18258 4868 18262 4924
rect 18262 4868 18318 4924
rect 18318 4868 18322 4924
rect 18258 4864 18322 4868
rect 18338 4924 18402 4928
rect 18338 4868 18342 4924
rect 18342 4868 18398 4924
rect 18398 4868 18402 4924
rect 18338 4864 18402 4868
rect 5850 4380 5914 4384
rect 5850 4324 5854 4380
rect 5854 4324 5910 4380
rect 5910 4324 5914 4380
rect 5850 4320 5914 4324
rect 5930 4380 5994 4384
rect 5930 4324 5934 4380
rect 5934 4324 5990 4380
rect 5990 4324 5994 4380
rect 5930 4320 5994 4324
rect 6010 4380 6074 4384
rect 6010 4324 6014 4380
rect 6014 4324 6070 4380
rect 6070 4324 6074 4380
rect 6010 4320 6074 4324
rect 6090 4380 6154 4384
rect 6090 4324 6094 4380
rect 6094 4324 6150 4380
rect 6150 4324 6154 4380
rect 6090 4320 6154 4324
rect 10749 4380 10813 4384
rect 10749 4324 10753 4380
rect 10753 4324 10809 4380
rect 10809 4324 10813 4380
rect 10749 4320 10813 4324
rect 10829 4380 10893 4384
rect 10829 4324 10833 4380
rect 10833 4324 10889 4380
rect 10889 4324 10893 4380
rect 10829 4320 10893 4324
rect 10909 4380 10973 4384
rect 10909 4324 10913 4380
rect 10913 4324 10969 4380
rect 10969 4324 10973 4380
rect 10909 4320 10973 4324
rect 10989 4380 11053 4384
rect 10989 4324 10993 4380
rect 10993 4324 11049 4380
rect 11049 4324 11053 4380
rect 10989 4320 11053 4324
rect 15648 4380 15712 4384
rect 15648 4324 15652 4380
rect 15652 4324 15708 4380
rect 15708 4324 15712 4380
rect 15648 4320 15712 4324
rect 15728 4380 15792 4384
rect 15728 4324 15732 4380
rect 15732 4324 15788 4380
rect 15788 4324 15792 4380
rect 15728 4320 15792 4324
rect 15808 4380 15872 4384
rect 15808 4324 15812 4380
rect 15812 4324 15868 4380
rect 15868 4324 15872 4380
rect 15808 4320 15872 4324
rect 15888 4380 15952 4384
rect 15888 4324 15892 4380
rect 15892 4324 15948 4380
rect 15948 4324 15952 4380
rect 15888 4320 15952 4324
rect 20547 4380 20611 4384
rect 20547 4324 20551 4380
rect 20551 4324 20607 4380
rect 20607 4324 20611 4380
rect 20547 4320 20611 4324
rect 20627 4380 20691 4384
rect 20627 4324 20631 4380
rect 20631 4324 20687 4380
rect 20687 4324 20691 4380
rect 20627 4320 20691 4324
rect 20707 4380 20771 4384
rect 20707 4324 20711 4380
rect 20711 4324 20767 4380
rect 20767 4324 20771 4380
rect 20707 4320 20771 4324
rect 20787 4380 20851 4384
rect 20787 4324 20791 4380
rect 20791 4324 20847 4380
rect 20847 4324 20851 4380
rect 20787 4320 20851 4324
rect 3401 3836 3465 3840
rect 3401 3780 3405 3836
rect 3405 3780 3461 3836
rect 3461 3780 3465 3836
rect 3401 3776 3465 3780
rect 3481 3836 3545 3840
rect 3481 3780 3485 3836
rect 3485 3780 3541 3836
rect 3541 3780 3545 3836
rect 3481 3776 3545 3780
rect 3561 3836 3625 3840
rect 3561 3780 3565 3836
rect 3565 3780 3621 3836
rect 3621 3780 3625 3836
rect 3561 3776 3625 3780
rect 3641 3836 3705 3840
rect 3641 3780 3645 3836
rect 3645 3780 3701 3836
rect 3701 3780 3705 3836
rect 3641 3776 3705 3780
rect 8300 3836 8364 3840
rect 8300 3780 8304 3836
rect 8304 3780 8360 3836
rect 8360 3780 8364 3836
rect 8300 3776 8364 3780
rect 8380 3836 8444 3840
rect 8380 3780 8384 3836
rect 8384 3780 8440 3836
rect 8440 3780 8444 3836
rect 8380 3776 8444 3780
rect 8460 3836 8524 3840
rect 8460 3780 8464 3836
rect 8464 3780 8520 3836
rect 8520 3780 8524 3836
rect 8460 3776 8524 3780
rect 8540 3836 8604 3840
rect 8540 3780 8544 3836
rect 8544 3780 8600 3836
rect 8600 3780 8604 3836
rect 8540 3776 8604 3780
rect 13199 3836 13263 3840
rect 13199 3780 13203 3836
rect 13203 3780 13259 3836
rect 13259 3780 13263 3836
rect 13199 3776 13263 3780
rect 13279 3836 13343 3840
rect 13279 3780 13283 3836
rect 13283 3780 13339 3836
rect 13339 3780 13343 3836
rect 13279 3776 13343 3780
rect 13359 3836 13423 3840
rect 13359 3780 13363 3836
rect 13363 3780 13419 3836
rect 13419 3780 13423 3836
rect 13359 3776 13423 3780
rect 13439 3836 13503 3840
rect 13439 3780 13443 3836
rect 13443 3780 13499 3836
rect 13499 3780 13503 3836
rect 13439 3776 13503 3780
rect 18098 3836 18162 3840
rect 18098 3780 18102 3836
rect 18102 3780 18158 3836
rect 18158 3780 18162 3836
rect 18098 3776 18162 3780
rect 18178 3836 18242 3840
rect 18178 3780 18182 3836
rect 18182 3780 18238 3836
rect 18238 3780 18242 3836
rect 18178 3776 18242 3780
rect 18258 3836 18322 3840
rect 18258 3780 18262 3836
rect 18262 3780 18318 3836
rect 18318 3780 18322 3836
rect 18258 3776 18322 3780
rect 18338 3836 18402 3840
rect 18338 3780 18342 3836
rect 18342 3780 18398 3836
rect 18398 3780 18402 3836
rect 18338 3776 18402 3780
rect 5850 3292 5914 3296
rect 5850 3236 5854 3292
rect 5854 3236 5910 3292
rect 5910 3236 5914 3292
rect 5850 3232 5914 3236
rect 5930 3292 5994 3296
rect 5930 3236 5934 3292
rect 5934 3236 5990 3292
rect 5990 3236 5994 3292
rect 5930 3232 5994 3236
rect 6010 3292 6074 3296
rect 6010 3236 6014 3292
rect 6014 3236 6070 3292
rect 6070 3236 6074 3292
rect 6010 3232 6074 3236
rect 6090 3292 6154 3296
rect 6090 3236 6094 3292
rect 6094 3236 6150 3292
rect 6150 3236 6154 3292
rect 6090 3232 6154 3236
rect 10749 3292 10813 3296
rect 10749 3236 10753 3292
rect 10753 3236 10809 3292
rect 10809 3236 10813 3292
rect 10749 3232 10813 3236
rect 10829 3292 10893 3296
rect 10829 3236 10833 3292
rect 10833 3236 10889 3292
rect 10889 3236 10893 3292
rect 10829 3232 10893 3236
rect 10909 3292 10973 3296
rect 10909 3236 10913 3292
rect 10913 3236 10969 3292
rect 10969 3236 10973 3292
rect 10909 3232 10973 3236
rect 10989 3292 11053 3296
rect 10989 3236 10993 3292
rect 10993 3236 11049 3292
rect 11049 3236 11053 3292
rect 10989 3232 11053 3236
rect 15648 3292 15712 3296
rect 15648 3236 15652 3292
rect 15652 3236 15708 3292
rect 15708 3236 15712 3292
rect 15648 3232 15712 3236
rect 15728 3292 15792 3296
rect 15728 3236 15732 3292
rect 15732 3236 15788 3292
rect 15788 3236 15792 3292
rect 15728 3232 15792 3236
rect 15808 3292 15872 3296
rect 15808 3236 15812 3292
rect 15812 3236 15868 3292
rect 15868 3236 15872 3292
rect 15808 3232 15872 3236
rect 15888 3292 15952 3296
rect 15888 3236 15892 3292
rect 15892 3236 15948 3292
rect 15948 3236 15952 3292
rect 15888 3232 15952 3236
rect 20547 3292 20611 3296
rect 20547 3236 20551 3292
rect 20551 3236 20607 3292
rect 20607 3236 20611 3292
rect 20547 3232 20611 3236
rect 20627 3292 20691 3296
rect 20627 3236 20631 3292
rect 20631 3236 20687 3292
rect 20687 3236 20691 3292
rect 20627 3232 20691 3236
rect 20707 3292 20771 3296
rect 20707 3236 20711 3292
rect 20711 3236 20767 3292
rect 20767 3236 20771 3292
rect 20707 3232 20771 3236
rect 20787 3292 20851 3296
rect 20787 3236 20791 3292
rect 20791 3236 20847 3292
rect 20847 3236 20851 3292
rect 20787 3232 20851 3236
rect 3401 2748 3465 2752
rect 3401 2692 3405 2748
rect 3405 2692 3461 2748
rect 3461 2692 3465 2748
rect 3401 2688 3465 2692
rect 3481 2748 3545 2752
rect 3481 2692 3485 2748
rect 3485 2692 3541 2748
rect 3541 2692 3545 2748
rect 3481 2688 3545 2692
rect 3561 2748 3625 2752
rect 3561 2692 3565 2748
rect 3565 2692 3621 2748
rect 3621 2692 3625 2748
rect 3561 2688 3625 2692
rect 3641 2748 3705 2752
rect 3641 2692 3645 2748
rect 3645 2692 3701 2748
rect 3701 2692 3705 2748
rect 3641 2688 3705 2692
rect 8300 2748 8364 2752
rect 8300 2692 8304 2748
rect 8304 2692 8360 2748
rect 8360 2692 8364 2748
rect 8300 2688 8364 2692
rect 8380 2748 8444 2752
rect 8380 2692 8384 2748
rect 8384 2692 8440 2748
rect 8440 2692 8444 2748
rect 8380 2688 8444 2692
rect 8460 2748 8524 2752
rect 8460 2692 8464 2748
rect 8464 2692 8520 2748
rect 8520 2692 8524 2748
rect 8460 2688 8524 2692
rect 8540 2748 8604 2752
rect 8540 2692 8544 2748
rect 8544 2692 8600 2748
rect 8600 2692 8604 2748
rect 8540 2688 8604 2692
rect 13199 2748 13263 2752
rect 13199 2692 13203 2748
rect 13203 2692 13259 2748
rect 13259 2692 13263 2748
rect 13199 2688 13263 2692
rect 13279 2748 13343 2752
rect 13279 2692 13283 2748
rect 13283 2692 13339 2748
rect 13339 2692 13343 2748
rect 13279 2688 13343 2692
rect 13359 2748 13423 2752
rect 13359 2692 13363 2748
rect 13363 2692 13419 2748
rect 13419 2692 13423 2748
rect 13359 2688 13423 2692
rect 13439 2748 13503 2752
rect 13439 2692 13443 2748
rect 13443 2692 13499 2748
rect 13499 2692 13503 2748
rect 13439 2688 13503 2692
rect 18098 2748 18162 2752
rect 18098 2692 18102 2748
rect 18102 2692 18158 2748
rect 18158 2692 18162 2748
rect 18098 2688 18162 2692
rect 18178 2748 18242 2752
rect 18178 2692 18182 2748
rect 18182 2692 18238 2748
rect 18238 2692 18242 2748
rect 18178 2688 18242 2692
rect 18258 2748 18322 2752
rect 18258 2692 18262 2748
rect 18262 2692 18318 2748
rect 18318 2692 18322 2748
rect 18258 2688 18322 2692
rect 18338 2748 18402 2752
rect 18338 2692 18342 2748
rect 18342 2692 18398 2748
rect 18398 2692 18402 2748
rect 18338 2688 18402 2692
rect 5850 2204 5914 2208
rect 5850 2148 5854 2204
rect 5854 2148 5910 2204
rect 5910 2148 5914 2204
rect 5850 2144 5914 2148
rect 5930 2204 5994 2208
rect 5930 2148 5934 2204
rect 5934 2148 5990 2204
rect 5990 2148 5994 2204
rect 5930 2144 5994 2148
rect 6010 2204 6074 2208
rect 6010 2148 6014 2204
rect 6014 2148 6070 2204
rect 6070 2148 6074 2204
rect 6010 2144 6074 2148
rect 6090 2204 6154 2208
rect 6090 2148 6094 2204
rect 6094 2148 6150 2204
rect 6150 2148 6154 2204
rect 6090 2144 6154 2148
rect 10749 2204 10813 2208
rect 10749 2148 10753 2204
rect 10753 2148 10809 2204
rect 10809 2148 10813 2204
rect 10749 2144 10813 2148
rect 10829 2204 10893 2208
rect 10829 2148 10833 2204
rect 10833 2148 10889 2204
rect 10889 2148 10893 2204
rect 10829 2144 10893 2148
rect 10909 2204 10973 2208
rect 10909 2148 10913 2204
rect 10913 2148 10969 2204
rect 10969 2148 10973 2204
rect 10909 2144 10973 2148
rect 10989 2204 11053 2208
rect 10989 2148 10993 2204
rect 10993 2148 11049 2204
rect 11049 2148 11053 2204
rect 10989 2144 11053 2148
rect 15648 2204 15712 2208
rect 15648 2148 15652 2204
rect 15652 2148 15708 2204
rect 15708 2148 15712 2204
rect 15648 2144 15712 2148
rect 15728 2204 15792 2208
rect 15728 2148 15732 2204
rect 15732 2148 15788 2204
rect 15788 2148 15792 2204
rect 15728 2144 15792 2148
rect 15808 2204 15872 2208
rect 15808 2148 15812 2204
rect 15812 2148 15868 2204
rect 15868 2148 15872 2204
rect 15808 2144 15872 2148
rect 15888 2204 15952 2208
rect 15888 2148 15892 2204
rect 15892 2148 15948 2204
rect 15948 2148 15952 2204
rect 15888 2144 15952 2148
rect 20547 2204 20611 2208
rect 20547 2148 20551 2204
rect 20551 2148 20607 2204
rect 20607 2148 20611 2204
rect 20547 2144 20611 2148
rect 20627 2204 20691 2208
rect 20627 2148 20631 2204
rect 20631 2148 20687 2204
rect 20687 2148 20691 2204
rect 20627 2144 20691 2148
rect 20707 2204 20771 2208
rect 20707 2148 20711 2204
rect 20711 2148 20767 2204
rect 20767 2148 20771 2204
rect 20707 2144 20771 2148
rect 20787 2204 20851 2208
rect 20787 2148 20791 2204
rect 20791 2148 20847 2204
rect 20847 2148 20851 2204
rect 20787 2144 20851 2148
<< metal4 >>
rect 3393 21248 3713 21808
rect 3393 21184 3401 21248
rect 3465 21184 3481 21248
rect 3545 21184 3561 21248
rect 3625 21184 3641 21248
rect 3705 21184 3713 21248
rect 3393 20160 3713 21184
rect 3393 20096 3401 20160
rect 3465 20096 3481 20160
rect 3545 20096 3561 20160
rect 3625 20096 3641 20160
rect 3705 20096 3713 20160
rect 3393 19072 3713 20096
rect 3393 19008 3401 19072
rect 3465 19008 3481 19072
rect 3545 19008 3561 19072
rect 3625 19008 3641 19072
rect 3705 19008 3713 19072
rect 3393 17984 3713 19008
rect 3393 17920 3401 17984
rect 3465 17920 3481 17984
rect 3545 17920 3561 17984
rect 3625 17920 3641 17984
rect 3705 17920 3713 17984
rect 3393 16896 3713 17920
rect 3393 16832 3401 16896
rect 3465 16832 3481 16896
rect 3545 16832 3561 16896
rect 3625 16832 3641 16896
rect 3705 16832 3713 16896
rect 3393 15808 3713 16832
rect 3393 15744 3401 15808
rect 3465 15744 3481 15808
rect 3545 15744 3561 15808
rect 3625 15744 3641 15808
rect 3705 15744 3713 15808
rect 3393 14720 3713 15744
rect 3393 14656 3401 14720
rect 3465 14656 3481 14720
rect 3545 14656 3561 14720
rect 3625 14656 3641 14720
rect 3705 14656 3713 14720
rect 3393 13632 3713 14656
rect 3393 13568 3401 13632
rect 3465 13568 3481 13632
rect 3545 13568 3561 13632
rect 3625 13568 3641 13632
rect 3705 13568 3713 13632
rect 3393 12544 3713 13568
rect 3393 12480 3401 12544
rect 3465 12480 3481 12544
rect 3545 12480 3561 12544
rect 3625 12480 3641 12544
rect 3705 12480 3713 12544
rect 3393 11456 3713 12480
rect 3393 11392 3401 11456
rect 3465 11392 3481 11456
rect 3545 11392 3561 11456
rect 3625 11392 3641 11456
rect 3705 11392 3713 11456
rect 3393 10368 3713 11392
rect 3393 10304 3401 10368
rect 3465 10304 3481 10368
rect 3545 10304 3561 10368
rect 3625 10304 3641 10368
rect 3705 10304 3713 10368
rect 3393 9280 3713 10304
rect 3393 9216 3401 9280
rect 3465 9216 3481 9280
rect 3545 9216 3561 9280
rect 3625 9216 3641 9280
rect 3705 9216 3713 9280
rect 3393 8192 3713 9216
rect 3393 8128 3401 8192
rect 3465 8128 3481 8192
rect 3545 8128 3561 8192
rect 3625 8128 3641 8192
rect 3705 8128 3713 8192
rect 3393 7104 3713 8128
rect 3393 7040 3401 7104
rect 3465 7040 3481 7104
rect 3545 7040 3561 7104
rect 3625 7040 3641 7104
rect 3705 7040 3713 7104
rect 3393 6016 3713 7040
rect 3393 5952 3401 6016
rect 3465 5952 3481 6016
rect 3545 5952 3561 6016
rect 3625 5952 3641 6016
rect 3705 5952 3713 6016
rect 3393 4928 3713 5952
rect 3393 4864 3401 4928
rect 3465 4864 3481 4928
rect 3545 4864 3561 4928
rect 3625 4864 3641 4928
rect 3705 4864 3713 4928
rect 3393 3840 3713 4864
rect 3393 3776 3401 3840
rect 3465 3776 3481 3840
rect 3545 3776 3561 3840
rect 3625 3776 3641 3840
rect 3705 3776 3713 3840
rect 3393 2752 3713 3776
rect 3393 2688 3401 2752
rect 3465 2688 3481 2752
rect 3545 2688 3561 2752
rect 3625 2688 3641 2752
rect 3705 2688 3713 2752
rect 3393 2128 3713 2688
rect 5842 21792 6162 21808
rect 5842 21728 5850 21792
rect 5914 21728 5930 21792
rect 5994 21728 6010 21792
rect 6074 21728 6090 21792
rect 6154 21728 6162 21792
rect 5842 20704 6162 21728
rect 5842 20640 5850 20704
rect 5914 20640 5930 20704
rect 5994 20640 6010 20704
rect 6074 20640 6090 20704
rect 6154 20640 6162 20704
rect 5842 19616 6162 20640
rect 5842 19552 5850 19616
rect 5914 19552 5930 19616
rect 5994 19552 6010 19616
rect 6074 19552 6090 19616
rect 6154 19552 6162 19616
rect 5842 18528 6162 19552
rect 5842 18464 5850 18528
rect 5914 18464 5930 18528
rect 5994 18464 6010 18528
rect 6074 18464 6090 18528
rect 6154 18464 6162 18528
rect 5842 17440 6162 18464
rect 5842 17376 5850 17440
rect 5914 17376 5930 17440
rect 5994 17376 6010 17440
rect 6074 17376 6090 17440
rect 6154 17376 6162 17440
rect 5842 16352 6162 17376
rect 5842 16288 5850 16352
rect 5914 16288 5930 16352
rect 5994 16288 6010 16352
rect 6074 16288 6090 16352
rect 6154 16288 6162 16352
rect 5842 15264 6162 16288
rect 5842 15200 5850 15264
rect 5914 15200 5930 15264
rect 5994 15200 6010 15264
rect 6074 15200 6090 15264
rect 6154 15200 6162 15264
rect 5842 14176 6162 15200
rect 5842 14112 5850 14176
rect 5914 14112 5930 14176
rect 5994 14112 6010 14176
rect 6074 14112 6090 14176
rect 6154 14112 6162 14176
rect 5842 13088 6162 14112
rect 5842 13024 5850 13088
rect 5914 13024 5930 13088
rect 5994 13024 6010 13088
rect 6074 13024 6090 13088
rect 6154 13024 6162 13088
rect 5842 12000 6162 13024
rect 5842 11936 5850 12000
rect 5914 11936 5930 12000
rect 5994 11936 6010 12000
rect 6074 11936 6090 12000
rect 6154 11936 6162 12000
rect 5842 10912 6162 11936
rect 5842 10848 5850 10912
rect 5914 10848 5930 10912
rect 5994 10848 6010 10912
rect 6074 10848 6090 10912
rect 6154 10848 6162 10912
rect 5842 9824 6162 10848
rect 5842 9760 5850 9824
rect 5914 9760 5930 9824
rect 5994 9760 6010 9824
rect 6074 9760 6090 9824
rect 6154 9760 6162 9824
rect 5842 8736 6162 9760
rect 5842 8672 5850 8736
rect 5914 8672 5930 8736
rect 5994 8672 6010 8736
rect 6074 8672 6090 8736
rect 6154 8672 6162 8736
rect 5842 7648 6162 8672
rect 5842 7584 5850 7648
rect 5914 7584 5930 7648
rect 5994 7584 6010 7648
rect 6074 7584 6090 7648
rect 6154 7584 6162 7648
rect 5842 6560 6162 7584
rect 5842 6496 5850 6560
rect 5914 6496 5930 6560
rect 5994 6496 6010 6560
rect 6074 6496 6090 6560
rect 6154 6496 6162 6560
rect 5842 5472 6162 6496
rect 5842 5408 5850 5472
rect 5914 5408 5930 5472
rect 5994 5408 6010 5472
rect 6074 5408 6090 5472
rect 6154 5408 6162 5472
rect 5842 4384 6162 5408
rect 5842 4320 5850 4384
rect 5914 4320 5930 4384
rect 5994 4320 6010 4384
rect 6074 4320 6090 4384
rect 6154 4320 6162 4384
rect 5842 3296 6162 4320
rect 5842 3232 5850 3296
rect 5914 3232 5930 3296
rect 5994 3232 6010 3296
rect 6074 3232 6090 3296
rect 6154 3232 6162 3296
rect 5842 2208 6162 3232
rect 5842 2144 5850 2208
rect 5914 2144 5930 2208
rect 5994 2144 6010 2208
rect 6074 2144 6090 2208
rect 6154 2144 6162 2208
rect 5842 2128 6162 2144
rect 8292 21248 8612 21808
rect 8292 21184 8300 21248
rect 8364 21184 8380 21248
rect 8444 21184 8460 21248
rect 8524 21184 8540 21248
rect 8604 21184 8612 21248
rect 8292 20160 8612 21184
rect 8292 20096 8300 20160
rect 8364 20096 8380 20160
rect 8444 20096 8460 20160
rect 8524 20096 8540 20160
rect 8604 20096 8612 20160
rect 8292 19072 8612 20096
rect 8292 19008 8300 19072
rect 8364 19008 8380 19072
rect 8444 19008 8460 19072
rect 8524 19008 8540 19072
rect 8604 19008 8612 19072
rect 8292 17984 8612 19008
rect 8292 17920 8300 17984
rect 8364 17920 8380 17984
rect 8444 17920 8460 17984
rect 8524 17920 8540 17984
rect 8604 17920 8612 17984
rect 8292 16896 8612 17920
rect 8292 16832 8300 16896
rect 8364 16832 8380 16896
rect 8444 16832 8460 16896
rect 8524 16832 8540 16896
rect 8604 16832 8612 16896
rect 8292 15808 8612 16832
rect 8292 15744 8300 15808
rect 8364 15744 8380 15808
rect 8444 15744 8460 15808
rect 8524 15744 8540 15808
rect 8604 15744 8612 15808
rect 8292 14720 8612 15744
rect 8292 14656 8300 14720
rect 8364 14656 8380 14720
rect 8444 14656 8460 14720
rect 8524 14656 8540 14720
rect 8604 14656 8612 14720
rect 8292 13632 8612 14656
rect 8292 13568 8300 13632
rect 8364 13568 8380 13632
rect 8444 13568 8460 13632
rect 8524 13568 8540 13632
rect 8604 13568 8612 13632
rect 8292 12544 8612 13568
rect 8292 12480 8300 12544
rect 8364 12480 8380 12544
rect 8444 12480 8460 12544
rect 8524 12480 8540 12544
rect 8604 12480 8612 12544
rect 8292 11456 8612 12480
rect 8292 11392 8300 11456
rect 8364 11392 8380 11456
rect 8444 11392 8460 11456
rect 8524 11392 8540 11456
rect 8604 11392 8612 11456
rect 8292 10368 8612 11392
rect 8292 10304 8300 10368
rect 8364 10304 8380 10368
rect 8444 10304 8460 10368
rect 8524 10304 8540 10368
rect 8604 10304 8612 10368
rect 8292 9280 8612 10304
rect 8292 9216 8300 9280
rect 8364 9216 8380 9280
rect 8444 9216 8460 9280
rect 8524 9216 8540 9280
rect 8604 9216 8612 9280
rect 8292 8192 8612 9216
rect 8292 8128 8300 8192
rect 8364 8128 8380 8192
rect 8444 8128 8460 8192
rect 8524 8128 8540 8192
rect 8604 8128 8612 8192
rect 8292 7104 8612 8128
rect 8292 7040 8300 7104
rect 8364 7040 8380 7104
rect 8444 7040 8460 7104
rect 8524 7040 8540 7104
rect 8604 7040 8612 7104
rect 8292 6016 8612 7040
rect 8292 5952 8300 6016
rect 8364 5952 8380 6016
rect 8444 5952 8460 6016
rect 8524 5952 8540 6016
rect 8604 5952 8612 6016
rect 8292 4928 8612 5952
rect 8292 4864 8300 4928
rect 8364 4864 8380 4928
rect 8444 4864 8460 4928
rect 8524 4864 8540 4928
rect 8604 4864 8612 4928
rect 8292 3840 8612 4864
rect 8292 3776 8300 3840
rect 8364 3776 8380 3840
rect 8444 3776 8460 3840
rect 8524 3776 8540 3840
rect 8604 3776 8612 3840
rect 8292 2752 8612 3776
rect 8292 2688 8300 2752
rect 8364 2688 8380 2752
rect 8444 2688 8460 2752
rect 8524 2688 8540 2752
rect 8604 2688 8612 2752
rect 8292 2128 8612 2688
rect 10741 21792 11061 21808
rect 10741 21728 10749 21792
rect 10813 21728 10829 21792
rect 10893 21728 10909 21792
rect 10973 21728 10989 21792
rect 11053 21728 11061 21792
rect 10741 20704 11061 21728
rect 10741 20640 10749 20704
rect 10813 20640 10829 20704
rect 10893 20640 10909 20704
rect 10973 20640 10989 20704
rect 11053 20640 11061 20704
rect 10741 19616 11061 20640
rect 10741 19552 10749 19616
rect 10813 19552 10829 19616
rect 10893 19552 10909 19616
rect 10973 19552 10989 19616
rect 11053 19552 11061 19616
rect 10741 18528 11061 19552
rect 10741 18464 10749 18528
rect 10813 18464 10829 18528
rect 10893 18464 10909 18528
rect 10973 18464 10989 18528
rect 11053 18464 11061 18528
rect 10741 17440 11061 18464
rect 10741 17376 10749 17440
rect 10813 17376 10829 17440
rect 10893 17376 10909 17440
rect 10973 17376 10989 17440
rect 11053 17376 11061 17440
rect 10741 16352 11061 17376
rect 10741 16288 10749 16352
rect 10813 16288 10829 16352
rect 10893 16288 10909 16352
rect 10973 16288 10989 16352
rect 11053 16288 11061 16352
rect 10741 15264 11061 16288
rect 10741 15200 10749 15264
rect 10813 15200 10829 15264
rect 10893 15200 10909 15264
rect 10973 15200 10989 15264
rect 11053 15200 11061 15264
rect 10741 14176 11061 15200
rect 10741 14112 10749 14176
rect 10813 14112 10829 14176
rect 10893 14112 10909 14176
rect 10973 14112 10989 14176
rect 11053 14112 11061 14176
rect 10741 13088 11061 14112
rect 10741 13024 10749 13088
rect 10813 13024 10829 13088
rect 10893 13024 10909 13088
rect 10973 13024 10989 13088
rect 11053 13024 11061 13088
rect 10741 12000 11061 13024
rect 10741 11936 10749 12000
rect 10813 11936 10829 12000
rect 10893 11936 10909 12000
rect 10973 11936 10989 12000
rect 11053 11936 11061 12000
rect 10741 10912 11061 11936
rect 10741 10848 10749 10912
rect 10813 10848 10829 10912
rect 10893 10848 10909 10912
rect 10973 10848 10989 10912
rect 11053 10848 11061 10912
rect 10741 9824 11061 10848
rect 10741 9760 10749 9824
rect 10813 9760 10829 9824
rect 10893 9760 10909 9824
rect 10973 9760 10989 9824
rect 11053 9760 11061 9824
rect 10741 8736 11061 9760
rect 10741 8672 10749 8736
rect 10813 8672 10829 8736
rect 10893 8672 10909 8736
rect 10973 8672 10989 8736
rect 11053 8672 11061 8736
rect 10741 7648 11061 8672
rect 10741 7584 10749 7648
rect 10813 7584 10829 7648
rect 10893 7584 10909 7648
rect 10973 7584 10989 7648
rect 11053 7584 11061 7648
rect 10741 6560 11061 7584
rect 10741 6496 10749 6560
rect 10813 6496 10829 6560
rect 10893 6496 10909 6560
rect 10973 6496 10989 6560
rect 11053 6496 11061 6560
rect 10741 5472 11061 6496
rect 10741 5408 10749 5472
rect 10813 5408 10829 5472
rect 10893 5408 10909 5472
rect 10973 5408 10989 5472
rect 11053 5408 11061 5472
rect 10741 4384 11061 5408
rect 10741 4320 10749 4384
rect 10813 4320 10829 4384
rect 10893 4320 10909 4384
rect 10973 4320 10989 4384
rect 11053 4320 11061 4384
rect 10741 3296 11061 4320
rect 10741 3232 10749 3296
rect 10813 3232 10829 3296
rect 10893 3232 10909 3296
rect 10973 3232 10989 3296
rect 11053 3232 11061 3296
rect 10741 2208 11061 3232
rect 10741 2144 10749 2208
rect 10813 2144 10829 2208
rect 10893 2144 10909 2208
rect 10973 2144 10989 2208
rect 11053 2144 11061 2208
rect 10741 2128 11061 2144
rect 13191 21248 13511 21808
rect 13191 21184 13199 21248
rect 13263 21184 13279 21248
rect 13343 21184 13359 21248
rect 13423 21184 13439 21248
rect 13503 21184 13511 21248
rect 13191 20160 13511 21184
rect 13191 20096 13199 20160
rect 13263 20096 13279 20160
rect 13343 20096 13359 20160
rect 13423 20096 13439 20160
rect 13503 20096 13511 20160
rect 13191 19072 13511 20096
rect 13191 19008 13199 19072
rect 13263 19008 13279 19072
rect 13343 19008 13359 19072
rect 13423 19008 13439 19072
rect 13503 19008 13511 19072
rect 13191 17984 13511 19008
rect 13191 17920 13199 17984
rect 13263 17920 13279 17984
rect 13343 17920 13359 17984
rect 13423 17920 13439 17984
rect 13503 17920 13511 17984
rect 13191 16896 13511 17920
rect 13191 16832 13199 16896
rect 13263 16832 13279 16896
rect 13343 16832 13359 16896
rect 13423 16832 13439 16896
rect 13503 16832 13511 16896
rect 13191 15808 13511 16832
rect 13191 15744 13199 15808
rect 13263 15744 13279 15808
rect 13343 15744 13359 15808
rect 13423 15744 13439 15808
rect 13503 15744 13511 15808
rect 13191 14720 13511 15744
rect 13191 14656 13199 14720
rect 13263 14656 13279 14720
rect 13343 14656 13359 14720
rect 13423 14656 13439 14720
rect 13503 14656 13511 14720
rect 13191 13632 13511 14656
rect 13191 13568 13199 13632
rect 13263 13568 13279 13632
rect 13343 13568 13359 13632
rect 13423 13568 13439 13632
rect 13503 13568 13511 13632
rect 13191 12544 13511 13568
rect 13191 12480 13199 12544
rect 13263 12480 13279 12544
rect 13343 12480 13359 12544
rect 13423 12480 13439 12544
rect 13503 12480 13511 12544
rect 13191 11456 13511 12480
rect 13191 11392 13199 11456
rect 13263 11392 13279 11456
rect 13343 11392 13359 11456
rect 13423 11392 13439 11456
rect 13503 11392 13511 11456
rect 13191 10368 13511 11392
rect 13191 10304 13199 10368
rect 13263 10304 13279 10368
rect 13343 10304 13359 10368
rect 13423 10304 13439 10368
rect 13503 10304 13511 10368
rect 13191 9280 13511 10304
rect 13191 9216 13199 9280
rect 13263 9216 13279 9280
rect 13343 9216 13359 9280
rect 13423 9216 13439 9280
rect 13503 9216 13511 9280
rect 13191 8192 13511 9216
rect 13191 8128 13199 8192
rect 13263 8128 13279 8192
rect 13343 8128 13359 8192
rect 13423 8128 13439 8192
rect 13503 8128 13511 8192
rect 13191 7104 13511 8128
rect 13191 7040 13199 7104
rect 13263 7040 13279 7104
rect 13343 7040 13359 7104
rect 13423 7040 13439 7104
rect 13503 7040 13511 7104
rect 13191 6016 13511 7040
rect 13191 5952 13199 6016
rect 13263 5952 13279 6016
rect 13343 5952 13359 6016
rect 13423 5952 13439 6016
rect 13503 5952 13511 6016
rect 13191 4928 13511 5952
rect 13191 4864 13199 4928
rect 13263 4864 13279 4928
rect 13343 4864 13359 4928
rect 13423 4864 13439 4928
rect 13503 4864 13511 4928
rect 13191 3840 13511 4864
rect 13191 3776 13199 3840
rect 13263 3776 13279 3840
rect 13343 3776 13359 3840
rect 13423 3776 13439 3840
rect 13503 3776 13511 3840
rect 13191 2752 13511 3776
rect 13191 2688 13199 2752
rect 13263 2688 13279 2752
rect 13343 2688 13359 2752
rect 13423 2688 13439 2752
rect 13503 2688 13511 2752
rect 13191 2128 13511 2688
rect 15640 21792 15960 21808
rect 15640 21728 15648 21792
rect 15712 21728 15728 21792
rect 15792 21728 15808 21792
rect 15872 21728 15888 21792
rect 15952 21728 15960 21792
rect 15640 20704 15960 21728
rect 15640 20640 15648 20704
rect 15712 20640 15728 20704
rect 15792 20640 15808 20704
rect 15872 20640 15888 20704
rect 15952 20640 15960 20704
rect 15640 19616 15960 20640
rect 15640 19552 15648 19616
rect 15712 19552 15728 19616
rect 15792 19552 15808 19616
rect 15872 19552 15888 19616
rect 15952 19552 15960 19616
rect 15640 18528 15960 19552
rect 15640 18464 15648 18528
rect 15712 18464 15728 18528
rect 15792 18464 15808 18528
rect 15872 18464 15888 18528
rect 15952 18464 15960 18528
rect 15640 17440 15960 18464
rect 15640 17376 15648 17440
rect 15712 17376 15728 17440
rect 15792 17376 15808 17440
rect 15872 17376 15888 17440
rect 15952 17376 15960 17440
rect 15640 16352 15960 17376
rect 15640 16288 15648 16352
rect 15712 16288 15728 16352
rect 15792 16288 15808 16352
rect 15872 16288 15888 16352
rect 15952 16288 15960 16352
rect 15640 15264 15960 16288
rect 15640 15200 15648 15264
rect 15712 15200 15728 15264
rect 15792 15200 15808 15264
rect 15872 15200 15888 15264
rect 15952 15200 15960 15264
rect 15640 14176 15960 15200
rect 15640 14112 15648 14176
rect 15712 14112 15728 14176
rect 15792 14112 15808 14176
rect 15872 14112 15888 14176
rect 15952 14112 15960 14176
rect 15640 13088 15960 14112
rect 15640 13024 15648 13088
rect 15712 13024 15728 13088
rect 15792 13024 15808 13088
rect 15872 13024 15888 13088
rect 15952 13024 15960 13088
rect 15640 12000 15960 13024
rect 15640 11936 15648 12000
rect 15712 11936 15728 12000
rect 15792 11936 15808 12000
rect 15872 11936 15888 12000
rect 15952 11936 15960 12000
rect 15640 10912 15960 11936
rect 15640 10848 15648 10912
rect 15712 10848 15728 10912
rect 15792 10848 15808 10912
rect 15872 10848 15888 10912
rect 15952 10848 15960 10912
rect 15640 9824 15960 10848
rect 15640 9760 15648 9824
rect 15712 9760 15728 9824
rect 15792 9760 15808 9824
rect 15872 9760 15888 9824
rect 15952 9760 15960 9824
rect 15640 8736 15960 9760
rect 15640 8672 15648 8736
rect 15712 8672 15728 8736
rect 15792 8672 15808 8736
rect 15872 8672 15888 8736
rect 15952 8672 15960 8736
rect 15640 7648 15960 8672
rect 15640 7584 15648 7648
rect 15712 7584 15728 7648
rect 15792 7584 15808 7648
rect 15872 7584 15888 7648
rect 15952 7584 15960 7648
rect 15640 6560 15960 7584
rect 15640 6496 15648 6560
rect 15712 6496 15728 6560
rect 15792 6496 15808 6560
rect 15872 6496 15888 6560
rect 15952 6496 15960 6560
rect 15640 5472 15960 6496
rect 15640 5408 15648 5472
rect 15712 5408 15728 5472
rect 15792 5408 15808 5472
rect 15872 5408 15888 5472
rect 15952 5408 15960 5472
rect 15640 4384 15960 5408
rect 15640 4320 15648 4384
rect 15712 4320 15728 4384
rect 15792 4320 15808 4384
rect 15872 4320 15888 4384
rect 15952 4320 15960 4384
rect 15640 3296 15960 4320
rect 15640 3232 15648 3296
rect 15712 3232 15728 3296
rect 15792 3232 15808 3296
rect 15872 3232 15888 3296
rect 15952 3232 15960 3296
rect 15640 2208 15960 3232
rect 15640 2144 15648 2208
rect 15712 2144 15728 2208
rect 15792 2144 15808 2208
rect 15872 2144 15888 2208
rect 15952 2144 15960 2208
rect 15640 2128 15960 2144
rect 18090 21248 18410 21808
rect 18090 21184 18098 21248
rect 18162 21184 18178 21248
rect 18242 21184 18258 21248
rect 18322 21184 18338 21248
rect 18402 21184 18410 21248
rect 18090 20160 18410 21184
rect 18090 20096 18098 20160
rect 18162 20096 18178 20160
rect 18242 20096 18258 20160
rect 18322 20096 18338 20160
rect 18402 20096 18410 20160
rect 18090 19072 18410 20096
rect 18090 19008 18098 19072
rect 18162 19008 18178 19072
rect 18242 19008 18258 19072
rect 18322 19008 18338 19072
rect 18402 19008 18410 19072
rect 18090 17984 18410 19008
rect 18090 17920 18098 17984
rect 18162 17920 18178 17984
rect 18242 17920 18258 17984
rect 18322 17920 18338 17984
rect 18402 17920 18410 17984
rect 18090 16896 18410 17920
rect 18090 16832 18098 16896
rect 18162 16832 18178 16896
rect 18242 16832 18258 16896
rect 18322 16832 18338 16896
rect 18402 16832 18410 16896
rect 18090 15808 18410 16832
rect 18090 15744 18098 15808
rect 18162 15744 18178 15808
rect 18242 15744 18258 15808
rect 18322 15744 18338 15808
rect 18402 15744 18410 15808
rect 18090 14720 18410 15744
rect 18090 14656 18098 14720
rect 18162 14656 18178 14720
rect 18242 14656 18258 14720
rect 18322 14656 18338 14720
rect 18402 14656 18410 14720
rect 18090 13632 18410 14656
rect 18090 13568 18098 13632
rect 18162 13568 18178 13632
rect 18242 13568 18258 13632
rect 18322 13568 18338 13632
rect 18402 13568 18410 13632
rect 18090 12544 18410 13568
rect 18090 12480 18098 12544
rect 18162 12480 18178 12544
rect 18242 12480 18258 12544
rect 18322 12480 18338 12544
rect 18402 12480 18410 12544
rect 18090 11456 18410 12480
rect 18090 11392 18098 11456
rect 18162 11392 18178 11456
rect 18242 11392 18258 11456
rect 18322 11392 18338 11456
rect 18402 11392 18410 11456
rect 18090 10368 18410 11392
rect 18090 10304 18098 10368
rect 18162 10304 18178 10368
rect 18242 10304 18258 10368
rect 18322 10304 18338 10368
rect 18402 10304 18410 10368
rect 18090 9280 18410 10304
rect 18090 9216 18098 9280
rect 18162 9216 18178 9280
rect 18242 9216 18258 9280
rect 18322 9216 18338 9280
rect 18402 9216 18410 9280
rect 18090 8192 18410 9216
rect 18090 8128 18098 8192
rect 18162 8128 18178 8192
rect 18242 8128 18258 8192
rect 18322 8128 18338 8192
rect 18402 8128 18410 8192
rect 18090 7104 18410 8128
rect 18090 7040 18098 7104
rect 18162 7040 18178 7104
rect 18242 7040 18258 7104
rect 18322 7040 18338 7104
rect 18402 7040 18410 7104
rect 18090 6016 18410 7040
rect 18090 5952 18098 6016
rect 18162 5952 18178 6016
rect 18242 5952 18258 6016
rect 18322 5952 18338 6016
rect 18402 5952 18410 6016
rect 18090 4928 18410 5952
rect 18090 4864 18098 4928
rect 18162 4864 18178 4928
rect 18242 4864 18258 4928
rect 18322 4864 18338 4928
rect 18402 4864 18410 4928
rect 18090 3840 18410 4864
rect 18090 3776 18098 3840
rect 18162 3776 18178 3840
rect 18242 3776 18258 3840
rect 18322 3776 18338 3840
rect 18402 3776 18410 3840
rect 18090 2752 18410 3776
rect 18090 2688 18098 2752
rect 18162 2688 18178 2752
rect 18242 2688 18258 2752
rect 18322 2688 18338 2752
rect 18402 2688 18410 2752
rect 18090 2128 18410 2688
rect 20539 21792 20859 21808
rect 20539 21728 20547 21792
rect 20611 21728 20627 21792
rect 20691 21728 20707 21792
rect 20771 21728 20787 21792
rect 20851 21728 20859 21792
rect 20539 20704 20859 21728
rect 20539 20640 20547 20704
rect 20611 20640 20627 20704
rect 20691 20640 20707 20704
rect 20771 20640 20787 20704
rect 20851 20640 20859 20704
rect 20539 19616 20859 20640
rect 20539 19552 20547 19616
rect 20611 19552 20627 19616
rect 20691 19552 20707 19616
rect 20771 19552 20787 19616
rect 20851 19552 20859 19616
rect 20539 18528 20859 19552
rect 20539 18464 20547 18528
rect 20611 18464 20627 18528
rect 20691 18464 20707 18528
rect 20771 18464 20787 18528
rect 20851 18464 20859 18528
rect 20539 17440 20859 18464
rect 20539 17376 20547 17440
rect 20611 17376 20627 17440
rect 20691 17376 20707 17440
rect 20771 17376 20787 17440
rect 20851 17376 20859 17440
rect 20539 16352 20859 17376
rect 20539 16288 20547 16352
rect 20611 16288 20627 16352
rect 20691 16288 20707 16352
rect 20771 16288 20787 16352
rect 20851 16288 20859 16352
rect 20539 15264 20859 16288
rect 20539 15200 20547 15264
rect 20611 15200 20627 15264
rect 20691 15200 20707 15264
rect 20771 15200 20787 15264
rect 20851 15200 20859 15264
rect 20539 14176 20859 15200
rect 20539 14112 20547 14176
rect 20611 14112 20627 14176
rect 20691 14112 20707 14176
rect 20771 14112 20787 14176
rect 20851 14112 20859 14176
rect 20539 13088 20859 14112
rect 20539 13024 20547 13088
rect 20611 13024 20627 13088
rect 20691 13024 20707 13088
rect 20771 13024 20787 13088
rect 20851 13024 20859 13088
rect 20539 12000 20859 13024
rect 20539 11936 20547 12000
rect 20611 11936 20627 12000
rect 20691 11936 20707 12000
rect 20771 11936 20787 12000
rect 20851 11936 20859 12000
rect 20539 10912 20859 11936
rect 20539 10848 20547 10912
rect 20611 10848 20627 10912
rect 20691 10848 20707 10912
rect 20771 10848 20787 10912
rect 20851 10848 20859 10912
rect 20539 9824 20859 10848
rect 20539 9760 20547 9824
rect 20611 9760 20627 9824
rect 20691 9760 20707 9824
rect 20771 9760 20787 9824
rect 20851 9760 20859 9824
rect 20539 8736 20859 9760
rect 20539 8672 20547 8736
rect 20611 8672 20627 8736
rect 20691 8672 20707 8736
rect 20771 8672 20787 8736
rect 20851 8672 20859 8736
rect 20539 7648 20859 8672
rect 20539 7584 20547 7648
rect 20611 7584 20627 7648
rect 20691 7584 20707 7648
rect 20771 7584 20787 7648
rect 20851 7584 20859 7648
rect 20539 6560 20859 7584
rect 20539 6496 20547 6560
rect 20611 6496 20627 6560
rect 20691 6496 20707 6560
rect 20771 6496 20787 6560
rect 20851 6496 20859 6560
rect 20539 5472 20859 6496
rect 20539 5408 20547 5472
rect 20611 5408 20627 5472
rect 20691 5408 20707 5472
rect 20771 5408 20787 5472
rect 20851 5408 20859 5472
rect 20539 4384 20859 5408
rect 20539 4320 20547 4384
rect 20611 4320 20627 4384
rect 20691 4320 20707 4384
rect 20771 4320 20787 4384
rect 20851 4320 20859 4384
rect 20539 3296 20859 4320
rect 20539 3232 20547 3296
rect 20611 3232 20627 3296
rect 20691 3232 20707 3296
rect 20771 3232 20787 3296
rect 20851 3232 20859 3296
rect 20539 2208 20859 3232
rect 20539 2144 20547 2208
rect 20611 2144 20627 2208
rect 20691 2144 20707 2208
rect 20771 2144 20787 2208
rect 20851 2144 20859 2208
rect 20539 2128 20859 2144
use sky130_fd_sc_hd__clkbuf_4  fanout52 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10672 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11408 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout54
timestamp 1704896540
transform 1 0 17664 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout55
timestamp 1704896540
transform 1 0 17756 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout56
timestamp 1704896540
transform 1 0 17204 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17572 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout58
timestamp 1704896540
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout59
timestamp 1704896540
transform -1 0 7636 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout60
timestamp 1704896540
transform 1 0 7636 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout61
timestamp 1704896540
transform -1 0 2944 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout62
timestamp 1704896540
transform -1 0 4508 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout63
timestamp 1704896540
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout64
timestamp 1704896540
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout65
timestamp 1704896540
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout66
timestamp 1704896540
transform -1 0 3680 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout67
timestamp 1704896540
transform -1 0 9476 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout68
timestamp 1704896540
transform -1 0 20240 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout69
timestamp 1704896540
transform 1 0 19872 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout70
timestamp 1704896540
transform -1 0 8004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout71
timestamp 1704896540
transform -1 0 13984 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2300 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_69
timestamp 1704896540
transform 1 0 7452 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_77
timestamp 1704896540
transform 1 0 8188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1704896540
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_106
timestamp 1704896540
transform 1 0 10856 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1704896540
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_113
timestamp 1704896540
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_125
timestamp 1704896540
transform 1 0 12604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_133
timestamp 1704896540
transform 1 0 13340 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1704896540
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_141
timestamp 1704896540
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_153
timestamp 1704896540
transform 1 0 15180 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_161
timestamp 1704896540
transform 1 0 15916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1704896540
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_169
timestamp 1704896540
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_181
timestamp 1704896540
transform 1 0 17756 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_189
timestamp 1704896540
transform 1 0 18492 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1704896540
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_197
timestamp 1704896540
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_44
timestamp 1704896540
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_57
timestamp 1704896540
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_80
timestamp 1704896540
transform 1 0 8464 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_88
timestamp 1704896540
transform 1 0 9200 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_110
timestamp 1704896540
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_139
timestamp 1704896540
transform 1 0 13892 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_151
timestamp 1704896540
transform 1 0 14996 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_163 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1704896540
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_169
timestamp 1704896540
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_194
timestamp 1704896540
transform 1 0 18952 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_23
timestamp 1704896540
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_62
timestamp 1704896540
transform 1 0 6808 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_70
timestamp 1704896540
transform 1 0 7544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_78
timestamp 1704896540
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_97
timestamp 1704896540
transform 1 0 10028 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_125
timestamp 1704896540
transform 1 0 12604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_137
timestamp 1704896540
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1704896540
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_153
timestamp 1704896540
transform 1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1704896540
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1704896540
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1704896540
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_197
timestamp 1704896540
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_205
timestamp 1704896540
transform 1 0 19964 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_69
timestamp 1704896540
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_73
timestamp 1704896540
transform 1 0 7820 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_82
timestamp 1704896540
transform 1 0 8648 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_94
timestamp 1704896540
transform 1 0 9752 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_106
timestamp 1704896540
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1704896540
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1704896540
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1704896540
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1704896540
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1704896540
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1704896540
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1704896540
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_181
timestamp 1704896540
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_189
timestamp 1704896540
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_32
timestamp 1704896540
transform 1 0 4048 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_37
timestamp 1704896540
transform 1 0 4508 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_48
timestamp 1704896540
transform 1 0 5520 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_60
timestamp 1704896540
transform 1 0 6624 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_66
timestamp 1704896540
transform 1 0 7176 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_80
timestamp 1704896540
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_97
timestamp 1704896540
transform 1 0 10028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_101
timestamp 1704896540
transform 1 0 10396 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_122
timestamp 1704896540
transform 1 0 12328 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_134
timestamp 1704896540
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_157
timestamp 1704896540
transform 1 0 15548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_169
timestamp 1704896540
transform 1 0 16652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_181
timestamp 1704896540
transform 1 0 17756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1704896540
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1704896540
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_209
timestamp 1704896540
transform 1 0 20332 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1704896540
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_78
timestamp 1704896540
transform 1 0 8280 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_90
timestamp 1704896540
transform 1 0 9384 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_95
timestamp 1704896540
transform 1 0 9844 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_107
timestamp 1704896540
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1704896540
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1704896540
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_125
timestamp 1704896540
transform 1 0 12604 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_133
timestamp 1704896540
transform 1 0 13340 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_152
timestamp 1704896540
transform 1 0 15088 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_209
timestamp 1704896540
transform 1 0 20332 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_15
timestamp 1704896540
transform 1 0 2484 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_23
timestamp 1704896540
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_45
timestamp 1704896540
transform 1 0 5244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_57
timestamp 1704896540
transform 1 0 6348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_69
timestamp 1704896540
transform 1 0 7452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_132
timestamp 1704896540
transform 1 0 13248 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_186
timestamp 1704896540
transform 1 0 18216 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_194
timestamp 1704896540
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_197
timestamp 1704896540
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_205
timestamp 1704896540
transform 1 0 19964 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_57
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_63
timestamp 1704896540
transform 1 0 6900 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_75
timestamp 1704896540
transform 1 0 8004 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_87
timestamp 1704896540
transform 1 0 9108 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1704896540
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1704896540
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1704896540
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1704896540
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1704896540
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1704896540
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1704896540
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1704896540
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1704896540
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_169
timestamp 1704896540
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_179
timestamp 1704896540
transform 1 0 17572 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_187
timestamp 1704896540
transform 1 0 18308 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_11
timestamp 1704896540
transform 1 0 2116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_20
timestamp 1704896540
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_37
timestamp 1704896540
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_97
timestamp 1704896540
transform 1 0 10028 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_108
timestamp 1704896540
transform 1 0 11040 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_120
timestamp 1704896540
transform 1 0 12144 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_132
timestamp 1704896540
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_141
timestamp 1704896540
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_147
timestamp 1704896540
transform 1 0 14628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_159
timestamp 1704896540
transform 1 0 15732 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_171
timestamp 1704896540
transform 1 0 16836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_183
timestamp 1704896540
transform 1 0 17940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1704896540
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_197
timestamp 1704896540
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_205
timestamp 1704896540
transform 1 0 19964 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_44
timestamp 1704896540
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_57
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_65
timestamp 1704896540
transform 1 0 7084 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1704896540
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_81
timestamp 1704896540
transform 1 0 8556 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1704896540
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_113
timestamp 1704896540
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_119
timestamp 1704896540
transform 1 0 12052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_124
timestamp 1704896540
transform 1 0 12512 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_129
timestamp 1704896540
transform 1 0 12972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_151
timestamp 1704896540
transform 1 0 14996 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_157
timestamp 1704896540
transform 1 0 15548 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_165
timestamp 1704896540
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_172
timestamp 1704896540
transform 1 0 16928 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_184
timestamp 1704896540
transform 1 0 18032 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_208
timestamp 1704896540
transform 1 0 20240 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_3
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_11
timestamp 1704896540
transform 1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_37
timestamp 1704896540
transform 1 0 4508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_47
timestamp 1704896540
transform 1 0 5428 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_55
timestamp 1704896540
transform 1 0 6164 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_80
timestamp 1704896540
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_91
timestamp 1704896540
transform 1 0 9476 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_96
timestamp 1704896540
transform 1 0 9936 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1704896540
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_141
timestamp 1704896540
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 1704896540
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1704896540
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_209
timestamp 1704896540
transform 1 0 20332 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1704896540
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1704896540
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1704896540
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1704896540
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1704896540
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_57
timestamp 1704896540
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_65
timestamp 1704896540
transform 1 0 7084 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_70
timestamp 1704896540
transform 1 0 7544 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_92
timestamp 1704896540
transform 1 0 9568 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_104
timestamp 1704896540
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_113
timestamp 1704896540
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_119
timestamp 1704896540
transform 1 0 12052 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_123
timestamp 1704896540
transform 1 0 12420 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_134
timestamp 1704896540
transform 1 0 13432 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_140
timestamp 1704896540
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_147
timestamp 1704896540
transform 1 0 14628 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_159
timestamp 1704896540
transform 1 0 15732 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_163
timestamp 1704896540
transform 1 0 16100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1704896540
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_169
timestamp 1704896540
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_178
timestamp 1704896540
transform 1 0 17480 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_188
timestamp 1704896540
transform 1 0 18400 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1704896540
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1704896540
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_50
timestamp 1704896540
transform 1 0 5704 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_58
timestamp 1704896540
transform 1 0 6440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_63
timestamp 1704896540
transform 1 0 6900 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_71
timestamp 1704896540
transform 1 0 7636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1704896540
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1704896540
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1704896540
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1704896540
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1704896540
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1704896540
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1704896540
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1704896540
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1704896540
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1704896540
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1704896540
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1704896540
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1704896540
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_197
timestamp 1704896540
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_205
timestamp 1704896540
transform 1 0 19964 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_25
timestamp 1704896540
transform 1 0 3404 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_33
timestamp 1704896540
transform 1 0 4140 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1704896540
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1704896540
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1704896540
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1704896540
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1704896540
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1704896540
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_113
timestamp 1704896540
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_121
timestamp 1704896540
transform 1 0 12236 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_126
timestamp 1704896540
transform 1 0 12696 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_130
timestamp 1704896540
transform 1 0 13064 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_134
timestamp 1704896540
transform 1 0 13432 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_146
timestamp 1704896540
transform 1 0 14536 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_158
timestamp 1704896540
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 1704896540
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1704896540
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1704896540
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1704896540
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_205
timestamp 1704896540
transform 1 0 19964 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_209
timestamp 1704896540
transform 1 0 20332 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1704896540
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_43
timestamp 1704896540
transform 1 0 5060 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_55
timestamp 1704896540
transform 1 0 6164 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_67
timestamp 1704896540
transform 1 0 7268 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_71
timestamp 1704896540
transform 1 0 7636 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_75
timestamp 1704896540
transform 1 0 8004 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1704896540
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_94
timestamp 1704896540
transform 1 0 9752 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_98
timestamp 1704896540
transform 1 0 10120 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_104
timestamp 1704896540
transform 1 0 10672 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_146
timestamp 1704896540
transform 1 0 14536 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_168
timestamp 1704896540
transform 1 0 16560 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_190
timestamp 1704896540
transform 1 0 18584 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_197
timestamp 1704896540
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_205
timestamp 1704896540
transform 1 0 19964 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_3
timestamp 1704896540
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_11
timestamp 1704896540
transform 1 0 2116 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1704896540
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1704896540
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1704896540
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1704896540
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1704896540
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_108
timestamp 1704896540
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_117
timestamp 1704896540
transform 1 0 11868 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_129
timestamp 1704896540
transform 1 0 12972 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_137
timestamp 1704896540
transform 1 0 13708 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_141
timestamp 1704896540
transform 1 0 14076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_153
timestamp 1704896540
transform 1 0 15180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_165
timestamp 1704896540
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_169
timestamp 1704896540
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_173
timestamp 1704896540
transform 1 0 17020 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1704896540
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_15
timestamp 1704896540
transform 1 0 2484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_20
timestamp 1704896540
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_41
timestamp 1704896540
transform 1 0 4876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_49
timestamp 1704896540
transform 1 0 5612 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_75
timestamp 1704896540
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1704896540
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_91
timestamp 1704896540
transform 1 0 9476 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_97
timestamp 1704896540
transform 1 0 10028 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_102
timestamp 1704896540
transform 1 0 10488 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_114
timestamp 1704896540
transform 1 0 11592 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_126
timestamp 1704896540
transform 1 0 12696 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_138
timestamp 1704896540
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_146
timestamp 1704896540
transform 1 0 14536 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_154
timestamp 1704896540
transform 1 0 15272 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_175
timestamp 1704896540
transform 1 0 17204 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_187
timestamp 1704896540
transform 1 0 18308 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1704896540
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1704896540
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_209
timestamp 1704896540
transform 1 0 20332 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_3
timestamp 1704896540
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_13
timestamp 1704896540
transform 1 0 2300 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_23
timestamp 1704896540
transform 1 0 3220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_29
timestamp 1704896540
transform 1 0 3772 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_34
timestamp 1704896540
transform 1 0 4232 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_46
timestamp 1704896540
transform 1 0 5336 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_52
timestamp 1704896540
transform 1 0 5888 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1704896540
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1704896540
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1704896540
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1704896540
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1704896540
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1704896540
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_113
timestamp 1704896540
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_120
timestamp 1704896540
transform 1 0 12144 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_128
timestamp 1704896540
transform 1 0 12880 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_151
timestamp 1704896540
transform 1 0 14996 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_163
timestamp 1704896540
transform 1 0 16100 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1704896540
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1704896540
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_181
timestamp 1704896540
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_189
timestamp 1704896540
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1704896540
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1704896540
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1704896540
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_43
timestamp 1704896540
transform 1 0 5060 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_58
timestamp 1704896540
transform 1 0 6440 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_70
timestamp 1704896540
transform 1 0 7544 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_82
timestamp 1704896540
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1704896540
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_109
timestamp 1704896540
transform 1 0 11132 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_135
timestamp 1704896540
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1704896540
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_141
timestamp 1704896540
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_167
timestamp 1704896540
transform 1 0 16468 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_191
timestamp 1704896540
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1704896540
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_197
timestamp 1704896540
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_205
timestamp 1704896540
transform 1 0 19964 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1704896540
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1704896540
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1704896540
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_45
timestamp 1704896540
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_53
timestamp 1704896540
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_57
timestamp 1704896540
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_61
timestamp 1704896540
transform 1 0 6716 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_65
timestamp 1704896540
transform 1 0 7084 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_76
timestamp 1704896540
transform 1 0 8096 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_104
timestamp 1704896540
transform 1 0 10672 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_108
timestamp 1704896540
transform 1 0 11040 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_113
timestamp 1704896540
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_122
timestamp 1704896540
transform 1 0 12328 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_134
timestamp 1704896540
transform 1 0 13432 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_146
timestamp 1704896540
transform 1 0 14536 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_158
timestamp 1704896540
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1704896540
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_189
timestamp 1704896540
transform 1 0 18492 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_201
timestamp 1704896540
transform 1 0 19596 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_209
timestamp 1704896540
transform 1 0 20332 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_3
timestamp 1704896540
transform 1 0 1380 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_16
timestamp 1704896540
transform 1 0 2576 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_41
timestamp 1704896540
transform 1 0 4876 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_45
timestamp 1704896540
transform 1 0 5244 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_50
timestamp 1704896540
transform 1 0 5704 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_62
timestamp 1704896540
transform 1 0 6808 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_74
timestamp 1704896540
transform 1 0 7912 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1704896540
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_85
timestamp 1704896540
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_131
timestamp 1704896540
transform 1 0 13156 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1704896540
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_161
timestamp 1704896540
transform 1 0 15916 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_173
timestamp 1704896540
transform 1 0 17020 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_187
timestamp 1704896540
transform 1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1704896540
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_197
timestamp 1704896540
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_205
timestamp 1704896540
transform 1 0 19964 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_6
timestamp 1704896540
transform 1 0 1656 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_32
timestamp 1704896540
transform 1 0 4048 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_44
timestamp 1704896540
transform 1 0 5152 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1704896540
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_69
timestamp 1704896540
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1704896540
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1704896540
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1704896540
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1704896540
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_125
timestamp 1704896540
transform 1 0 12604 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_131
timestamp 1704896540
transform 1 0 13156 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_135
timestamp 1704896540
transform 1 0 13524 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_144
timestamp 1704896540
transform 1 0 14352 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_156
timestamp 1704896540
transform 1 0 15456 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1704896540
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_181
timestamp 1704896540
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_189
timestamp 1704896540
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1704896540
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1704896540
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1704896540
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1704896540
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_41
timestamp 1704896540
transform 1 0 4876 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_45
timestamp 1704896540
transform 1 0 5244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_57
timestamp 1704896540
transform 1 0 6348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_69
timestamp 1704896540
transform 1 0 7452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 1704896540
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1704896540
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1704896540
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1704896540
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1704896540
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1704896540
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1704896540
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_161
timestamp 1704896540
transform 1 0 15916 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1704896540
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1704896540
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1704896540
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_209
timestamp 1704896540
transform 1 0 20332 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_3
timestamp 1704896540
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_7
timestamp 1704896540
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_11
timestamp 1704896540
transform 1 0 2116 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_19
timestamp 1704896540
transform 1 0 2852 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_42
timestamp 1704896540
transform 1 0 4968 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_50
timestamp 1704896540
transform 1 0 5704 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_80
timestamp 1704896540
transform 1 0 8464 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_85
timestamp 1704896540
transform 1 0 8924 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_89
timestamp 1704896540
transform 1 0 9292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_110
timestamp 1704896540
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_120
timestamp 1704896540
transform 1 0 12144 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_128
timestamp 1704896540
transform 1 0 12880 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1704896540
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1704896540
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1704896540
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_169
timestamp 1704896540
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_173
timestamp 1704896540
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_32
timestamp 1704896540
transform 1 0 4048 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_40
timestamp 1704896540
transform 1 0 4784 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_75
timestamp 1704896540
transform 1 0 8004 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 1704896540
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_105
timestamp 1704896540
transform 1 0 10764 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp 1704896540
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_144
timestamp 1704896540
transform 1 0 14352 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_190
timestamp 1704896540
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_197
timestamp 1704896540
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1704896540
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1704896540
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1704896540
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1704896540
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_51
timestamp 1704896540
transform 1 0 5796 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1704896540
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_57
timestamp 1704896540
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_62
timestamp 1704896540
transform 1 0 6808 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_85
timestamp 1704896540
transform 1 0 8924 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_96
timestamp 1704896540
transform 1 0 9936 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_108
timestamp 1704896540
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_113
timestamp 1704896540
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_119
timestamp 1704896540
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_123
timestamp 1704896540
transform 1 0 12420 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_135
timestamp 1704896540
transform 1 0 13524 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_147
timestamp 1704896540
transform 1 0 14628 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_159
timestamp 1704896540
transform 1 0 15732 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1704896540
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1704896540
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_181
timestamp 1704896540
transform 1 0 17756 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_209
timestamp 1704896540
transform 1 0 20332 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1704896540
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_15
timestamp 1704896540
transform 1 0 2484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_19
timestamp 1704896540
transform 1 0 2852 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_25
timestamp 1704896540
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_29
timestamp 1704896540
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_33
timestamp 1704896540
transform 1 0 4140 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_37
timestamp 1704896540
transform 1 0 4508 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_43
timestamp 1704896540
transform 1 0 5060 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_55
timestamp 1704896540
transform 1 0 6164 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_67
timestamp 1704896540
transform 1 0 7268 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_78
timestamp 1704896540
transform 1 0 8280 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1704896540
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_97
timestamp 1704896540
transform 1 0 10028 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_106
timestamp 1704896540
transform 1 0 10856 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_118
timestamp 1704896540
transform 1 0 11960 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_130
timestamp 1704896540
transform 1 0 13064 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1704896540
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1704896540
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_153
timestamp 1704896540
transform 1 0 15180 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_178
timestamp 1704896540
transform 1 0 17480 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_190
timestamp 1704896540
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_197
timestamp 1704896540
transform 1 0 19228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_201
timestamp 1704896540
transform 1 0 19596 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_208
timestamp 1704896540
transform 1 0 20240 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_3
timestamp 1704896540
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_7
timestamp 1704896540
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_11
timestamp 1704896540
transform 1 0 2116 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_19
timestamp 1704896540
transform 1 0 2852 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1704896540
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1704896540
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1704896540
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1704896540
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1704896540
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_69
timestamp 1704896540
transform 1 0 7452 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_75
timestamp 1704896540
transform 1 0 8004 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_100
timestamp 1704896540
transform 1 0 10304 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_106
timestamp 1704896540
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_117
timestamp 1704896540
transform 1 0 11868 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_129
timestamp 1704896540
transform 1 0 12972 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_135
timestamp 1704896540
transform 1 0 13524 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_139
timestamp 1704896540
transform 1 0 13892 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_151
timestamp 1704896540
transform 1 0 14996 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_159
timestamp 1704896540
transform 1 0 15732 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_163
timestamp 1704896540
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1704896540
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_169
timestamp 1704896540
transform 1 0 16652 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_173
timestamp 1704896540
transform 1 0 17020 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_185
timestamp 1704896540
transform 1 0 18124 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_189
timestamp 1704896540
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_3
timestamp 1704896540
transform 1 0 1380 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1704896540
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1704896540
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_53
timestamp 1704896540
transform 1 0 5980 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_74
timestamp 1704896540
transform 1 0 7912 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_82
timestamp 1704896540
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1704896540
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1704896540
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_109
timestamp 1704896540
transform 1 0 11132 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_161
timestamp 1704896540
transform 1 0 15916 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_173
timestamp 1704896540
transform 1 0 17020 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_185
timestamp 1704896540
transform 1 0 18124 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1704896540
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1704896540
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_205
timestamp 1704896540
transform 1 0 19964 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1704896540
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1704896540
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_27
timestamp 1704896540
transform 1 0 3588 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_31
timestamp 1704896540
transform 1 0 3956 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_52
timestamp 1704896540
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_57
timestamp 1704896540
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_63
timestamp 1704896540
transform 1 0 6900 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_84
timestamp 1704896540
transform 1 0 8832 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_88
timestamp 1704896540
transform 1 0 9200 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_109
timestamp 1704896540
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1704896540
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1704896540
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_137
timestamp 1704896540
transform 1 0 13708 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_143
timestamp 1704896540
transform 1 0 14260 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_147
timestamp 1704896540
transform 1 0 14628 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_163
timestamp 1704896540
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1704896540
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1704896540
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_181
timestamp 1704896540
transform 1 0 17756 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_202
timestamp 1704896540
transform 1 0 19688 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_3
timestamp 1704896540
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_7
timestamp 1704896540
transform 1 0 1748 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_11
timestamp 1704896540
transform 1 0 2116 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_23
timestamp 1704896540
transform 1 0 3220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1704896540
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1704896540
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_41
timestamp 1704896540
transform 1 0 4876 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_64
timestamp 1704896540
transform 1 0 6992 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_76
timestamp 1704896540
transform 1 0 8096 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1704896540
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_97
timestamp 1704896540
transform 1 0 10028 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_120
timestamp 1704896540
transform 1 0 12144 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_132
timestamp 1704896540
transform 1 0 13248 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1704896540
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1704896540
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_165
timestamp 1704896540
transform 1 0 16284 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_170
timestamp 1704896540
transform 1 0 16744 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_176
timestamp 1704896540
transform 1 0 17296 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_182
timestamp 1704896540
transform 1 0 17848 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1704896540
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_197
timestamp 1704896540
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_205
timestamp 1704896540
transform 1 0 19964 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_23
timestamp 1704896540
transform 1 0 3220 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_46
timestamp 1704896540
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_54
timestamp 1704896540
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1704896540
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_69
timestamp 1704896540
transform 1 0 7452 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_97
timestamp 1704896540
transform 1 0 10028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_109
timestamp 1704896540
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_133
timestamp 1704896540
transform 1 0 13340 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_145
timestamp 1704896540
transform 1 0 14444 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_157
timestamp 1704896540
transform 1 0 15548 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_165
timestamp 1704896540
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1704896540
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_181
timestamp 1704896540
transform 1 0 17756 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_203
timestamp 1704896540
transform 1 0 19780 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_209
timestamp 1704896540
transform 1 0 20332 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1704896540
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1704896540
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1704896540
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_29
timestamp 1704896540
transform 1 0 3772 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_33
timestamp 1704896540
transform 1 0 4140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_45
timestamp 1704896540
transform 1 0 5244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_57
timestamp 1704896540
transform 1 0 6348 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_80
timestamp 1704896540
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_88
timestamp 1704896540
transform 1 0 9200 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_100
timestamp 1704896540
transform 1 0 10304 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_112
timestamp 1704896540
transform 1 0 11408 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1704896540
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_153
timestamp 1704896540
transform 1 0 15180 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_178
timestamp 1704896540
transform 1 0 17480 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_187
timestamp 1704896540
transform 1 0 18308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1704896540
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_197
timestamp 1704896540
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_205
timestamp 1704896540
transform 1 0 19964 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1704896540
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1704896540
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_47
timestamp 1704896540
transform 1 0 5428 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1704896540
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_57
timestamp 1704896540
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_65
timestamp 1704896540
transform 1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1704896540
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1704896540
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_125
timestamp 1704896540
transform 1 0 12604 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_129
timestamp 1704896540
transform 1 0 12972 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_150
timestamp 1704896540
transform 1 0 14904 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_162
timestamp 1704896540
transform 1 0 16008 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1704896540
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_181
timestamp 1704896540
transform 1 0 17756 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_7
timestamp 1704896540
transform 1 0 1748 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_19
timestamp 1704896540
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1704896540
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_41
timestamp 1704896540
transform 1 0 4876 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_47
timestamp 1704896540
transform 1 0 5428 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_68
timestamp 1704896540
transform 1 0 7360 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_75
timestamp 1704896540
transform 1 0 8004 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1704896540
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_94
timestamp 1704896540
transform 1 0 9752 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_126
timestamp 1704896540
transform 1 0 12696 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_134
timestamp 1704896540
transform 1 0 13432 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_161
timestamp 1704896540
transform 1 0 15916 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_169
timestamp 1704896540
transform 1 0 16652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_194
timestamp 1704896540
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_197
timestamp 1704896540
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1704896540
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_27
timestamp 1704896540
transform 1 0 3588 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_35
timestamp 1704896540
transform 1 0 4324 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_43
timestamp 1704896540
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1704896540
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_63
timestamp 1704896540
transform 1 0 6900 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_71
timestamp 1704896540
transform 1 0 7636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_83
timestamp 1704896540
transform 1 0 8740 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_91
timestamp 1704896540
transform 1 0 9476 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_99
timestamp 1704896540
transform 1 0 10212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1704896540
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_119
timestamp 1704896540
transform 1 0 12052 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_127
timestamp 1704896540
transform 1 0 12788 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_139
timestamp 1704896540
transform 1 0 13892 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_147
timestamp 1704896540
transform 1 0 14628 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_155
timestamp 1704896540
transform 1 0 15364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1704896540
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_175
timestamp 1704896540
transform 1 0 17204 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_183
timestamp 1704896540
transform 1 0 17940 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_195
timestamp 1704896540
transform 1 0 19044 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_203
timestamp 1704896540
transform 1 0 19780 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 20148 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1704896540
transform -1 0 19872 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1704896540
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1704896540
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1704896540
transform 1 0 20056 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1704896540
transform 1 0 20056 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1704896540
transform -1 0 20424 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1704896540
transform -1 0 19872 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1704896540
transform -1 0 20424 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1704896540
transform -1 0 20424 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1704896540
transform -1 0 20424 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1704896540
transform -1 0 20424 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1704896540
transform -1 0 20424 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1704896540
transform 1 0 20056 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1704896540
transform 1 0 20056 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1704896540
transform -1 0 19044 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1704896540
transform 1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1704896540
transform -1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1704896540
transform -1 0 11316 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1704896540
transform -1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1704896540
transform 1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1704896540
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1704896540
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1704896540
transform -1 0 20424 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1704896540
transform 1 0 19504 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1704896540
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1704896540
transform -1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1704896540
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1704896540
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1704896540
transform 1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1704896540
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output33
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 1704896540
transform 1 0 19228 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1704896540
transform 1 0 17388 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1704896540
transform -1 0 12788 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1704896540
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1704896540
transform -1 0 10212 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1704896540
transform -1 0 5060 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1704896540
transform 1 0 3772 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1704896540
transform -1 0 2484 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output42
timestamp 1704896540
transform -1 0 20424 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output43
timestamp 1704896540
transform 1 0 19872 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output44
timestamp 1704896540
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output45
timestamp 1704896540
transform 1 0 14812 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output46
timestamp 1704896540
transform 1 0 14076 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output47
timestamp 1704896540
transform 1 0 8924 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output48
timestamp 1704896540
transform 1 0 7084 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output49
timestamp 1704896540
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output50
timestamp 1704896540
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1704896540
transform -1 0 1748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_36
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_37
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 20700 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_38
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 20700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_39
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 20700 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_40
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 20700 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_41
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 20700 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_42
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 20700 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_43
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 20700 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_44
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 20700 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_45
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 20700 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_46
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 20700 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_47
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 20700 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_48
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 20700 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_49
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 20700 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_50
timestamp 1704896540
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 20700 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_51
timestamp 1704896540
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 20700 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_52
timestamp 1704896540
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 20700 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_53
timestamp 1704896540
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 20700 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_54
timestamp 1704896540
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 20700 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_55
timestamp 1704896540
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 20700 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_56
timestamp 1704896540
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 20700 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_57
timestamp 1704896540
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 20700 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_58
timestamp 1704896540
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 20700 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_59
timestamp 1704896540
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 20700 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_60
timestamp 1704896540
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 20700 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_61
timestamp 1704896540
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 20700 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_62
timestamp 1704896540
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 20700 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_63
timestamp 1704896540
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 20700 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_64
timestamp 1704896540
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1704896540
transform -1 0 20700 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_65
timestamp 1704896540
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1704896540
transform -1 0 20700 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_66
timestamp 1704896540
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1704896540
transform -1 0 20700 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_67
timestamp 1704896540
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1704896540
transform -1 0 20700 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_68
timestamp 1704896540
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1704896540
transform -1 0 20700 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_69
timestamp 1704896540
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1704896540
transform -1 0 20700 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_70
timestamp 1704896540
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1704896540
transform -1 0 20700 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_71
timestamp 1704896540
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1704896540
transform -1 0 20700 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_75
timestamp 1704896540
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_76
timestamp 1704896540
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_77
timestamp 1704896540
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 1704896540
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_79
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_80
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_81
timestamp 1704896540
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_82
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_83
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_84
timestamp 1704896540
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_85
timestamp 1704896540
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_86
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_87
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_88
timestamp 1704896540
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_89
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_90
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_91
timestamp 1704896540
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_92
timestamp 1704896540
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_93
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_94
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_95
timestamp 1704896540
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_96
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_97
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_98
timestamp 1704896540
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_99
timestamp 1704896540
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_100
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_101
timestamp 1704896540
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_102
timestamp 1704896540
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_103
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_104
timestamp 1704896540
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_105
timestamp 1704896540
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_106
timestamp 1704896540
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_107
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_108
timestamp 1704896540
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_109
timestamp 1704896540
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_110
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_111
timestamp 1704896540
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_112
timestamp 1704896540
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_113
timestamp 1704896540
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_114
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_115
timestamp 1704896540
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_116
timestamp 1704896540
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_117
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_118
timestamp 1704896540
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_119
timestamp 1704896540
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_120
timestamp 1704896540
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_121
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_122
timestamp 1704896540
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_123
timestamp 1704896540
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_124
timestamp 1704896540
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_125
timestamp 1704896540
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_126
timestamp 1704896540
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_127
timestamp 1704896540
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_128
timestamp 1704896540
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_129
timestamp 1704896540
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_130
timestamp 1704896540
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_131
timestamp 1704896540
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_132
timestamp 1704896540
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_133
timestamp 1704896540
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_134
timestamp 1704896540
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_135
timestamp 1704896540
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_136
timestamp 1704896540
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_137
timestamp 1704896540
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_138
timestamp 1704896540
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_139
timestamp 1704896540
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_140
timestamp 1704896540
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_141
timestamp 1704896540
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_142
timestamp 1704896540
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_143
timestamp 1704896540
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_144
timestamp 1704896540
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_145
timestamp 1704896540
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_146
timestamp 1704896540
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_147
timestamp 1704896540
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_148
timestamp 1704896540
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_149
timestamp 1704896540
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_150
timestamp 1704896540
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_151
timestamp 1704896540
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_152
timestamp 1704896540
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_153
timestamp 1704896540
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_154
timestamp 1704896540
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_155
timestamp 1704896540
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_156
timestamp 1704896540
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_157
timestamp 1704896540
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_158
timestamp 1704896540
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_159
timestamp 1704896540
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_160
timestamp 1704896540
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_161
timestamp 1704896540
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_162
timestamp 1704896540
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_163
timestamp 1704896540
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_164
timestamp 1704896540
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_165
timestamp 1704896540
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_166
timestamp 1704896540
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_167
timestamp 1704896540
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_168
timestamp 1704896540
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_169
timestamp 1704896540
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_170
timestamp 1704896540
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_171
timestamp 1704896540
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_172
timestamp 1704896540
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_173
timestamp 1704896540
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_174
timestamp 1704896540
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_175
timestamp 1704896540
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_176
timestamp 1704896540
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_177
timestamp 1704896540
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_178
timestamp 1704896540
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_179
timestamp 1704896540
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_180
timestamp 1704896540
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_181
timestamp 1704896540
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_182
timestamp 1704896540
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_183
timestamp 1704896540
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_184
timestamp 1704896540
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_185
timestamp 1704896540
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_186
timestamp 1704896540
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_187
timestamp 1704896540
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_188
timestamp 1704896540
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_189
timestamp 1704896540
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_190
timestamp 1704896540
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_191
timestamp 1704896540
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_192
timestamp 1704896540
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_193
timestamp 1704896540
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_194
timestamp 1704896540
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_195
timestamp 1704896540
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_196
timestamp 1704896540
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_197
timestamp 1704896540
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_198
timestamp 1704896540
transform 1 0 3680 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_199
timestamp 1704896540
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_200
timestamp 1704896540
transform 1 0 8832 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_201
timestamp 1704896540
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_202
timestamp 1704896540
transform 1 0 13984 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_203
timestamp 1704896540
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_204
timestamp 1704896540
transform 1 0 19136 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fa_1  x1_x1_x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17112 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  x1_x1_x2
timestamp 1704896540
transform 1 0 17020 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  x1_x1_x3
timestamp 1704896540
transform 1 0 17204 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  x1_x1_x4
timestamp 1704896540
transform 1 0 17112 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  x1_x1_x5
timestamp 1704896540
transform 1 0 17112 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  x1_x1_x6
timestamp 1704896540
transform 1 0 14076 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  x1_x1_x7
timestamp 1704896540
transform 1 0 13616 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  x1_x1_x8
timestamp 1704896540
transform 1 0 14076 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  x1_x1_x9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18584 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x1_x10
timestamp 1704896540
transform 1 0 18584 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x1_x11
timestamp 1704896540
transform 1 0 18584 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x1_x12
timestamp 1704896540
transform 1 0 18584 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x1_x13
timestamp 1704896540
transform 1 0 18584 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x1_x14
timestamp 1704896540
transform 1 0 18584 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x1_x15
timestamp 1704896540
transform 1 0 16652 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x1_x16
timestamp 1704896540
transform 1 0 18492 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x1_x17
timestamp 1704896540
transform 1 0 18584 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_1  x1_x1_x29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 19688 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x1_x1_x110
timestamp 1704896540
transform 1 0 18492 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x1
timestamp 1704896540
transform 1 0 18584 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x2
timestamp 1704896540
transform 1 0 17848 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x3
timestamp 1704896540
transform 1 0 17940 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  x1_x2_x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17020 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  x1_x2_x5
timestamp 1704896540
transform 1 0 15456 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  x1_x2_x6
timestamp 1704896540
transform 1 0 15548 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  x1_x2_x7
timestamp 1704896540
transform 1 0 17020 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  x1_x2_x8
timestamp 1704896540
transform 1 0 10672 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  x1_x2_x9
timestamp 1704896540
transform 1 0 18308 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x1_x2_x10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 19228 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x1_x2_x11
timestamp 1704896540
transform 1 0 18216 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x1_x2_x12
timestamp 1704896540
transform 1 0 18032 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x1_x2_x13
timestamp 1704896540
transform 1 0 17388 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x1_x2_x14
timestamp 1704896540
transform 1 0 16468 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x1_x2_x15
timestamp 1704896540
transform 1 0 16744 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  x1_x2_x16_x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17664 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x1_x2_x16_x9
timestamp 1704896540
transform 1 0 17204 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x1_x2_x16_x10
timestamp 1704896540
transform -1 0 17664 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  x1_x2_x17_x1
timestamp 1704896540
transform 1 0 15640 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x1_x2_x17_x9
timestamp 1704896540
transform 1 0 14904 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x1_x2_x17_x10
timestamp 1704896540
transform 1 0 15180 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x1_x2_x18
timestamp 1704896540
transform 1 0 15272 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x19
timestamp 1704896540
transform 1 0 14076 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_1  x1_x2_x20
timestamp 1704896540
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x1_x2_x21
timestamp 1704896540
transform 1 0 13892 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x22
timestamp 1704896540
transform 1 0 14076 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x23
timestamp 1704896540
transform 1 0 13156 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x24
timestamp 1704896540
transform 1 0 12972 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x25
timestamp 1704896540
transform 1 0 11684 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x26
timestamp 1704896540
transform 1 0 11592 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  x1_x2_x27
timestamp 1704896540
transform 1 0 10764 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  x1_x2_x28
timestamp 1704896540
transform 1 0 9292 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  x1_x2_x29
timestamp 1704896540
transform 1 0 13248 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x1_x2_x30
timestamp 1704896540
transform -1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x1_x2_x31
timestamp 1704896540
transform 1 0 14076 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x1_x2_x32
timestamp 1704896540
transform 1 0 13800 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x1_x2_x33
timestamp 1704896540
transform 1 0 11316 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x1_x2_x34
timestamp 1704896540
transform 1 0 10488 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  x1_x2_x35_x1
timestamp 1704896540
transform 1 0 14076 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x1_x2_x35_x9
timestamp 1704896540
transform 1 0 13156 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x1_x2_x35_x10
timestamp 1704896540
transform -1 0 13708 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  x1_x2_x36_x1
timestamp 1704896540
transform 1 0 10580 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x1_x2_x36_x9
timestamp 1704896540
transform -1 0 10120 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x1_x2_x36_x10
timestamp 1704896540
transform -1 0 10028 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x1_x2_x37
timestamp 1704896540
transform 1 0 11684 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x1_x2_x38
timestamp 1704896540
transform 1 0 11040 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  x1_x2_x39_x1
timestamp 1704896540
transform 1 0 7912 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x1_x2_x39_x9
timestamp 1704896540
transform -1 0 8464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x1_x2_x39_x10
timestamp 1704896540
transform -1 0 8188 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__dfstp_1  x1_x2_x40
timestamp 1704896540
transform 1 0 9200 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  x1_x2_x41
timestamp 1704896540
transform 1 0 8924 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  x1_x2_x42
timestamp 1704896540
transform -1 0 9752 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  x1_x2_x43
timestamp 1704896540
transform 1 0 8372 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  x1_x2_x44
timestamp 1704896540
transform 1 0 2852 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  x1_x2_x45
timestamp 1704896540
transform 1 0 8096 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x46
timestamp 1704896540
transform 1 0 6624 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_1  x1_x2_x47
timestamp 1704896540
transform 1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x1_x2_x48
timestamp 1704896540
transform -1 0 8280 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x49
timestamp 1704896540
transform 1 0 6716 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x50
timestamp 1704896540
transform 1 0 4968 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x51
timestamp 1704896540
transform 1 0 4416 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x52
timestamp 1704896540
transform 1 0 4048 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x53
timestamp 1704896540
transform 1 0 3864 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  x1_x2_x54
timestamp 1704896540
transform 1 0 3036 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  x1_x2_x55
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  x1_x2_x56
timestamp 1704896540
transform -1 0 8648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x1_x2_x57
timestamp 1704896540
transform -1 0 5060 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x1_x2_x58
timestamp 1704896540
transform 1 0 5152 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x1_x2_x59
timestamp 1704896540
transform -1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x1_x2_x60
timestamp 1704896540
transform -1 0 4784 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x1_x2_x61
timestamp 1704896540
transform -1 0 4048 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  x1_x2_x62_x1
timestamp 1704896540
transform 1 0 4784 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x1_x2_x62_x9
timestamp 1704896540
transform -1 0 5244 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x1_x2_x62_x10
timestamp 1704896540
transform -1 0 4968 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  x1_x2_x63_x1
timestamp 1704896540
transform 1 0 4048 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x1_x2_x63_x9
timestamp 1704896540
transform -1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x1_x2_x63_x10
timestamp 1704896540
transform -1 0 3680 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x1_x2_x64
timestamp 1704896540
transform -1 0 5152 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x1_x2_x65
timestamp 1704896540
transform -1 0 5428 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  x1_x2_x67
timestamp 1704896540
transform 1 0 1472 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  x1_x2_x68
timestamp 1704896540
transform -1 0 3312 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  x1_x2_x69
timestamp 1704896540
transform -1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  x1_x2_x70
timestamp 1704896540
transform 1 0 1380 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x71
timestamp 1704896540
transform 1 0 16744 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_1  x1_x2_x72
timestamp 1704896540
transform -1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x73
timestamp 1704896540
transform -1 0 3220 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_1  x1_x2_x74
timestamp 1704896540
transform 1 0 1840 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x75
timestamp 1704896540
transform -1 0 3220 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  x1_x2_x76
timestamp 1704896540
transform -1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x2_x77
timestamp 1704896540
transform -1 0 17020 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x78
timestamp 1704896540
transform 1 0 15364 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__xor2_1  x1_x2_x79 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15088 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  x1_x2_x80
timestamp 1704896540
transform -1 0 14628 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x2_x81
timestamp 1704896540
transform -1 0 13892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x82
timestamp 1704896540
transform 1 0 14076 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__xor2_1  x1_x2_x83
timestamp 1704896540
transform 1 0 13340 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  x1_x2_x84
timestamp 1704896540
transform -1 0 12052 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x2_x85
timestamp 1704896540
transform -1 0 11408 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x86
timestamp 1704896540
transform 1 0 11408 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__xor2_1  x1_x2_x87
timestamp 1704896540
transform 1 0 10028 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  x1_x2_x88
timestamp 1704896540
transform -1 0 13984 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x2_x89
timestamp 1704896540
transform -1 0 12696 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x90
timestamp 1704896540
transform 1 0 8740 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__xor2_1  x1_x2_x91
timestamp 1704896540
transform 1 0 10764 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  x1_x2_x92
timestamp 1704896540
transform -1 0 9476 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x2_x93
timestamp 1704896540
transform -1 0 8740 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x94
timestamp 1704896540
transform 1 0 6440 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__xor2_1  x1_x2_x95
timestamp 1704896540
transform -1 0 9752 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  x1_x2_x96
timestamp 1704896540
transform -1 0 7728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x2_x97
timestamp 1704896540
transform -1 0 7176 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x98
timestamp 1704896540
transform 1 0 3312 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__xor2_1  x1_x2_x99
timestamp 1704896540
transform 1 0 5612 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  x1_x2_x100
timestamp 1704896540
transform -1 0 4508 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x2_x101
timestamp 1704896540
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x102
timestamp 1704896540
transform 1 0 3312 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__xor2_1  x1_x2_x103
timestamp 1704896540
transform 1 0 2576 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  x1_x2_x104
timestamp 1704896540
transform -1 0 3220 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x2_x105
timestamp 1704896540
transform -1 0 2576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x106
timestamp 1704896540
transform 1 0 14904 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__xor2_1  x1_x2_x107
timestamp 1704896540
transform 1 0 2300 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_4  x1_x2_x108 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14352 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x109
timestamp 1704896540
transform 1 0 16652 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x110
timestamp 1704896540
transform 1 0 15364 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  x1_x2_x111
timestamp 1704896540
transform 1 0 11224 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x112
timestamp 1704896540
transform 1 0 14720 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  x1_x2_x113
timestamp 1704896540
transform -1 0 6716 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x114
timestamp 1704896540
transform 1 0 9200 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x115
timestamp 1704896540
transform 1 0 10488 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x116
timestamp 1704896540
transform 1 0 11408 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x117
timestamp 1704896540
transform 1 0 12052 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x118
timestamp 1704896540
transform 1 0 15824 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__and2_0  x1_x2_x119_x1
timestamp 1704896540
transform 1 0 12696 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x1_x2_x119_x9
timestamp 1704896540
transform 1 0 12052 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x1_x2_x119_x10
timestamp 1704896540
transform -1 0 12696 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x120
timestamp 1704896540
transform 1 0 18584 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2_x121
timestamp 1704896540
transform 1 0 10396 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x3_x1
timestamp 1704896540
transform 1 0 3588 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x3_x2
timestamp 1704896540
transform -1 0 5336 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x3_x3
timestamp 1704896540
transform 1 0 4048 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x3_x4
timestamp 1704896540
transform 1 0 5152 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x3_x5
timestamp 1704896540
transform 1 0 6072 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x3_x6
timestamp 1704896540
transform 1 0 6992 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x3_x7
timestamp 1704896540
transform 1 0 8188 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x3_x8
timestamp 1704896540
transform 1 0 9292 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x3_x9
timestamp 1704896540
transform 1 0 10304 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x3_x10
timestamp 1704896540
transform -1 0 7360 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x3_x11
timestamp 1704896540
transform 1 0 11500 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x3_x12
timestamp 1704896540
transform 1 0 12144 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x3_x13
timestamp 1704896540
transform 1 0 13064 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x3_x14
timestamp 1704896540
transform 1 0 14076 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x3_x15
timestamp 1704896540
transform -1 0 8464 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x3_x16
timestamp 1704896540
transform 1 0 7360 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  x1_x3_x17
timestamp 1704896540
transform 1 0 4600 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x3_x18
timestamp 1704896540
transform -1 0 4140 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  x1_x3_x19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4600 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  x1_x3_x20
timestamp 1704896540
transform -1 0 9200 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x3_x21
timestamp 1704896540
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x3_x22
timestamp 1704896540
transform 1 0 3312 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x1_x3_x23
timestamp 1704896540
transform -1 0 3312 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x1_x3_x24
timestamp 1704896540
transform -1 0 3404 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  x1_x3_x25
timestamp 1704896540
transform 1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x3_x26
timestamp 1704896540
transform 1 0 2208 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  x1_x3_x27
timestamp 1704896540
transform -1 0 2484 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_16  x1_x3_x28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3404 0 -1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__dfrtp_1  x1_x4_x1
timestamp 1704896540
transform 1 0 7084 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x4_x2
timestamp 1704896540
transform 1 0 8924 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x4_x3
timestamp 1704896540
transform 1 0 9384 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x4_x4
timestamp 1704896540
transform 1 0 7820 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x4_x5
timestamp 1704896540
transform 1 0 8188 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x4_x6
timestamp 1704896540
transform 1 0 6164 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x4_x7
timestamp 1704896540
transform 1 0 6348 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x4_x8
timestamp 1704896540
transform 1 0 6624 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x4_x9
timestamp 1704896540
transform 1 0 6348 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x4_x10
timestamp 1704896540
transform 1 0 7728 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x4_x11
timestamp 1704896540
transform 1 0 9108 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x4_x12
timestamp 1704896540
transform 1 0 10120 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x4_x13
timestamp 1704896540
transform 1 0 11960 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x4_x14
timestamp 1704896540
transform 1 0 13156 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x4_x15
timestamp 1704896540
transform 1 0 14444 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x4_x16
timestamp 1704896540
transform 1 0 16284 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x17
timestamp 1704896540
transform -1 0 5244 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x18
timestamp 1704896540
transform -1 0 6164 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x19
timestamp 1704896540
transform -1 0 6808 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x20
timestamp 1704896540
transform -1 0 8648 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x21
timestamp 1704896540
transform -1 0 8924 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x22
timestamp 1704896540
transform -1 0 8464 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x23
timestamp 1704896540
transform -1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x24
timestamp 1704896540
transform -1 0 8096 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x25
timestamp 1704896540
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x26
timestamp 1704896540
transform -1 0 6256 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x27
timestamp 1704896540
transform -1 0 6164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x28
timestamp 1704896540
transform -1 0 6624 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x29
timestamp 1704896540
transform -1 0 7544 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x30
timestamp 1704896540
transform -1 0 9200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x31
timestamp 1704896540
transform -1 0 9936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x32
timestamp 1704896540
transform 1 0 12144 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x33
timestamp 1704896540
transform -1 0 12972 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x34
timestamp 1704896540
transform -1 0 14352 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x35
timestamp 1704896540
transform -1 0 14628 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x36
timestamp 1704896540
transform -1 0 7636 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x37
timestamp 1704896540
transform 1 0 6164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x38
timestamp 1704896540
transform 1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x39
timestamp 1704896540
transform -1 0 9476 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x40
timestamp 1704896540
transform -1 0 12512 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x41
timestamp 1704896540
transform -1 0 13432 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x1_x4_x42
timestamp 1704896540
transform 1 0 6808 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  x1_x4_x43
timestamp 1704896540
transform 1 0 6992 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x44
timestamp 1704896540
transform -1 0 8280 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  x1_x4_x45
timestamp 1704896540
transform 1 0 10488 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x46
timestamp 1704896540
transform -1 0 9936 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x1_x4_x47
timestamp 1704896540
transform 1 0 10580 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x48
timestamp 1704896540
transform -1 0 11316 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x1_x4_x49
timestamp 1704896540
transform 1 0 12144 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x50
timestamp 1704896540
transform 1 0 11868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  x1_x4_x51
timestamp 1704896540
transform -1 0 11868 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x52
timestamp 1704896540
transform -1 0 9752 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x1_x4_x53
timestamp 1704896540
transform 1 0 9752 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x54
timestamp 1704896540
transform -1 0 10488 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x1_x4_x55
timestamp 1704896540
transform 1 0 11316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x56
timestamp 1704896540
transform -1 0 8004 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x1_x4_x57
timestamp 1704896540
transform 1 0 8188 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x58
timestamp 1704896540
transform 1 0 7360 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  x1_x4_x59
timestamp 1704896540
transform -1 0 6900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x60
timestamp 1704896540
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x1_x4_x61
timestamp 1704896540
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x62
timestamp 1704896540
transform -1 0 9660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x1_x4_x63
timestamp 1704896540
transform 1 0 9568 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x64
timestamp 1704896540
transform 1 0 10948 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x1_x4_x65
timestamp 1704896540
transform -1 0 11040 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x66
timestamp 1704896540
transform 1 0 11776 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  x1_x4_x67
timestamp 1704896540
transform 1 0 11684 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x68
timestamp 1704896540
transform -1 0 14628 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x69
timestamp 1704896540
transform -1 0 15824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x70
timestamp 1704896540
transform -1 0 15548 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x1_x4_x71
timestamp 1704896540
transform 1 0 15824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x72
timestamp 1704896540
transform -1 0 16928 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x73
timestamp 1704896540
transform -1 0 17480 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x74
timestamp 1704896540
transform -1 0 17204 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x4_x75
timestamp 1704896540
transform 1 0 17756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x1_x4_x76
timestamp 1704896540
transform 1 0 4600 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x1_x4_x77
timestamp 1704896540
transform 1 0 4232 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_16  x1_x4_x78
timestamp 1704896540
transform 1 0 5060 0 1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_1  x1_x5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17112 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__buf_16  x1_x6
timestamp 1704896540
transform 1 0 2024 0 -1 14144
box -38 -48 2062 592
use sky130_fd_sc_hd__clkbuf_1  x1_x7
timestamp 1704896540
transform -1 0 18400 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x8
timestamp 1704896540
transform -1 0 1748 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  x1_x9
timestamp 1704896540
transform 1 0 1748 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  x1_x12
timestamp 1704896540
transform 1 0 18124 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  x1_x24
timestamp 1704896540
transform 1 0 17664 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_16  x1_x78
timestamp 1704896540
transform 1 0 18216 0 -1 7616
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_1  x2_x1
timestamp 1704896540
transform 1 0 1656 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  x2_x2
timestamp 1704896540
transform 1 0 2668 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x2_x3
timestamp 1704896540
transform -1 0 2668 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x2_x4
timestamp 1704896540
transform -1 0 3220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x2_x5
timestamp 1704896540
transform -1 0 3772 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x2_x6
timestamp 1704896540
transform -1 0 4232 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x2_x7
timestamp 1704896540
transform 1 0 4784 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x2_x8
timestamp 1704896540
transform -1 0 4784 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x2_x9
timestamp 1704896540
transform 1 0 4968 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x2_x10
timestamp 1704896540
transform -1 0 4968 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x2_x11
timestamp 1704896540
transform -1 0 5704 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x2_x12
timestamp 1704896540
transform -1 0 5244 0 1 13056
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 GND
port 0 nsew signal bidirectional
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 VDD
port 1 nsew signal bidirectional
flabel metal4 s 5842 2128 6162 21808 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 10741 2128 11061 21808 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 15640 2128 15960 21808 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 20539 2128 20859 21808 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 3393 2128 3713 21808 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 8292 2128 8612 21808 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 13191 2128 13511 21808 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 18090 2128 18410 21808 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal3 s 21080 19864 21880 19984 0 FreeSans 480 0 0 0 clk
port 4 nsew signal input
flabel metal3 s 21080 21496 21880 21616 0 FreeSans 480 0 0 0 clr
port 5 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 comp_clk
port 6 nsew signal output
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 comp_n
port 7 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 comp_p
port 8 nsew signal input
flabel metal3 s 21080 18232 21880 18352 0 FreeSans 480 0 0 0 done
port 9 nsew signal output
flabel metal3 s 21080 16600 21880 16720 0 FreeSans 480 0 0 0 obit1
port 10 nsew signal output
flabel metal3 s 21080 1912 21880 2032 0 FreeSans 480 0 0 0 obit10
port 11 nsew signal output
flabel metal3 s 21080 14968 21880 15088 0 FreeSans 480 0 0 0 obit2
port 12 nsew signal output
flabel metal3 s 21080 13336 21880 13456 0 FreeSans 480 0 0 0 obit3
port 13 nsew signal output
flabel metal3 s 21080 11704 21880 11824 0 FreeSans 480 0 0 0 obit4
port 14 nsew signal output
flabel metal3 s 21080 10072 21880 10192 0 FreeSans 480 0 0 0 obit5
port 15 nsew signal output
flabel metal3 s 21080 8440 21880 8560 0 FreeSans 480 0 0 0 obit6
port 16 nsew signal output
flabel metal3 s 21080 6808 21880 6928 0 FreeSans 480 0 0 0 obit7
port 17 nsew signal output
flabel metal3 s 21080 5176 21880 5296 0 FreeSans 480 0 0 0 obit8
port 18 nsew signal output
flabel metal3 s 21080 3544 21880 3664 0 FreeSans 480 0 0 0 obit9
port 19 nsew signal output
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 sw_n1
port 20 nsew signal output
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 sw_n2
port 21 nsew signal output
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 sw_n3
port 22 nsew signal output
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 sw_n4
port 23 nsew signal output
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 sw_n5
port 24 nsew signal output
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 sw_n6
port 25 nsew signal output
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 sw_n7
port 26 nsew signal output
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 sw_n8
port 27 nsew signal output
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 sw_n_sp1
port 28 nsew signal output
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 sw_n_sp2
port 29 nsew signal output
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 sw_n_sp3
port 30 nsew signal output
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 sw_n_sp4
port 31 nsew signal output
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 sw_n_sp5
port 32 nsew signal output
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 sw_n_sp6
port 33 nsew signal output
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 sw_n_sp7
port 34 nsew signal output
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 sw_n_sp8
port 35 nsew signal output
flabel metal2 s 570 0 626 800 0 FreeSans 224 90 0 0 sw_n_sp9
port 36 nsew signal output
flabel metal2 s 18602 23224 18658 24024 0 FreeSans 224 90 0 0 sw_p1
port 37 nsew signal output
flabel metal2 s 17314 23224 17370 24024 0 FreeSans 224 90 0 0 sw_p2
port 38 nsew signal output
flabel metal2 s 12162 23224 12218 24024 0 FreeSans 224 90 0 0 sw_p3
port 39 nsew signal output
flabel metal2 s 10874 23224 10930 24024 0 FreeSans 224 90 0 0 sw_p4
port 40 nsew signal output
flabel metal2 s 9586 23224 9642 24024 0 FreeSans 224 90 0 0 sw_p5
port 41 nsew signal output
flabel metal2 s 4434 23224 4490 24024 0 FreeSans 224 90 0 0 sw_p6
port 42 nsew signal output
flabel metal2 s 3146 23224 3202 24024 0 FreeSans 224 90 0 0 sw_p7
port 43 nsew signal output
flabel metal2 s 1858 23224 1914 24024 0 FreeSans 224 90 0 0 sw_p8
port 44 nsew signal output
flabel metal2 s 21178 23224 21234 24024 0 FreeSans 224 90 0 0 sw_p_sp1
port 45 nsew signal output
flabel metal2 s 19890 23224 19946 24024 0 FreeSans 224 90 0 0 sw_p_sp2
port 46 nsew signal output
flabel metal2 s 16026 23224 16082 24024 0 FreeSans 224 90 0 0 sw_p_sp3
port 47 nsew signal output
flabel metal2 s 14738 23224 14794 24024 0 FreeSans 224 90 0 0 sw_p_sp4
port 48 nsew signal output
flabel metal2 s 13450 23224 13506 24024 0 FreeSans 224 90 0 0 sw_p_sp5
port 49 nsew signal output
flabel metal2 s 8298 23224 8354 24024 0 FreeSans 224 90 0 0 sw_p_sp6
port 50 nsew signal output
flabel metal2 s 7010 23224 7066 24024 0 FreeSans 224 90 0 0 sw_p_sp7
port 51 nsew signal output
flabel metal2 s 5722 23224 5778 24024 0 FreeSans 224 90 0 0 sw_p_sp8
port 52 nsew signal output
flabel metal2 s 570 23224 626 24024 0 FreeSans 224 90 0 0 sw_p_sp9
port 53 nsew signal output
flabel metal3 s 0 21224 800 21344 0 FreeSans 480 0 0 0 sw_sample
port 54 nsew signal output
rlabel via1 10981 21760 10981 21760 0 VGND
rlabel metal1 10902 21216 10902 21216 0 VPWR
rlabel metal3 1579 6052 1579 6052 0 VDD
rlabel metal2 20378 19873 20378 19873 0 clk
rlabel metal2 19642 21233 19642 21233 0 clr
rlabel metal3 1096 2244 1096 2244 0 comp_clk
rlabel metal3 751 9860 751 9860 0 comp_n
rlabel metal3 1050 13668 1050 13668 0 comp_p
rlabel metal1 6900 12818 6900 12818 0 controller_clk
rlabel metal2 20286 18445 20286 18445 0 done
rlabel metal1 18078 19720 18078 19720 0 net1
rlabel metal2 20378 13498 20378 13498 0 net10
rlabel metal2 20378 12036 20378 12036 0 net11
rlabel metal2 20378 10234 20378 10234 0 net12
rlabel metal2 20378 8772 20378 8772 0 net13
rlabel metal2 20378 6596 20378 6596 0 net14
rlabel metal2 18446 5508 18446 5508 0 net15
rlabel metal2 20102 4250 20102 4250 0 net16
rlabel metal2 18998 2618 18998 2618 0 net17
rlabel metal2 17434 2890 17434 2890 0 net18
rlabel metal2 12558 2890 12558 2890 0 net19
rlabel metal1 19642 20774 19642 20774 0 net2
rlabel metal1 11201 2822 11201 2822 0 net20
rlabel metal1 10557 2618 10557 2618 0 net21
rlabel metal1 4761 3026 4761 3026 0 net22
rlabel via1 3243 4998 3243 4998 0 net23
rlabel metal1 1725 7174 1725 7174 0 net24
rlabel metal1 20378 2414 20378 2414 0 net25
rlabel metal1 19596 18054 19596 18054 0 net26
rlabel metal2 16100 9996 16100 9996 0 net27
rlabel metal1 15088 2414 15088 2414 0 net28
rlabel metal2 13570 4657 13570 4657 0 net29
rlabel metal2 1794 10948 1794 10948 0 net3
rlabel metal1 8556 2414 8556 2414 0 net30
rlabel metal1 6946 3366 6946 3366 0 net31
rlabel metal1 5888 2414 5888 2414 0 net32
rlabel metal1 1472 2414 1472 2414 0 net33
rlabel metal1 19113 21114 19113 21114 0 net34
rlabel metal1 17457 20026 17457 20026 0 net35
rlabel via1 12627 21114 12627 21114 0 net36
rlabel metal1 11339 20570 11339 20570 0 net37
rlabel metal1 10143 17306 10143 17306 0 net38
rlabel via1 4899 15130 4899 15130 0 net39
rlabel metal2 1518 12512 1518 12512 0 net4
rlabel metal1 3565 17850 3565 17850 0 net40
rlabel metal1 3151 15674 3151 15674 0 net41
rlabel metal1 20332 20570 20332 20570 0 net42
rlabel metal2 19734 20502 19734 20502 0 net43
rlabel metal2 16790 19041 16790 19041 0 net44
rlabel metal1 14996 21522 14996 21522 0 net45
rlabel metal1 13800 15674 13800 15674 0 net46
rlabel metal2 8832 19380 8832 19380 0 net47
rlabel metal1 6716 9486 6716 9486 0 net48
rlabel metal1 6072 21522 6072 21522 0 net49
rlabel metal2 1702 6256 1702 6256 0 net5
rlabel metal1 1472 19482 1472 19482 0 net50
rlabel metal1 2231 20910 2231 20910 0 net51
rlabel metal1 2622 7480 2622 7480 0 net52
rlabel metal1 10449 2346 10449 2346 0 net53
rlabel metal1 17710 3128 17710 3128 0 net54
rlabel metal1 19458 17680 19458 17680 0 net55
rlabel metal2 2162 18462 2162 18462 0 net56
rlabel metal1 17572 6086 17572 6086 0 net57
rlabel metal1 18584 6290 18584 6290 0 net58
rlabel metal1 7590 15334 7590 15334 0 net59
rlabel metal1 19987 17850 19987 17850 0 net6
rlabel metal1 16698 7752 16698 7752 0 net60
rlabel metal1 4370 2312 4370 2312 0 net61
rlabel metal1 9430 2482 9430 2482 0 net62
rlabel metal1 15962 3570 15962 3570 0 net63
rlabel metal1 16790 12716 16790 12716 0 net64
rlabel metal1 18814 17102 18814 17102 0 net65
rlabel via1 1965 18734 1965 18734 0 net66
rlabel metal1 8977 20502 8977 20502 0 net67
rlabel metal1 18446 16694 18446 16694 0 net68
rlabel metal1 18676 6834 18676 6834 0 net69
rlabel metal1 20194 16218 20194 16218 0 net7
rlabel metal2 4094 17918 4094 17918 0 net70
rlabel metal1 13386 20842 13386 20842 0 net71
rlabel metal2 20378 3468 20378 3468 0 net8
rlabel metal1 20102 15130 20102 15130 0 net9
rlabel metal2 20286 17085 20286 17085 0 obit1
rlabel metal2 20194 2397 20194 2397 0 obit10
rlabel metal1 19458 15334 19458 15334 0 obit2
rlabel via2 20194 13413 20194 13413 0 obit3
rlabel metal2 20194 11917 20194 11917 0 obit4
rlabel via2 20194 10149 20194 10149 0 obit5
rlabel metal2 20194 8653 20194 8653 0 obit6
rlabel metal2 20194 6749 20194 6749 0 obit7
rlabel metal2 20286 5389 20286 5389 0 obit8
rlabel via2 20286 3621 20286 3621 0 obit9
rlabel metal2 18630 1520 18630 1520 0 sw_n1
rlabel metal2 17342 1520 17342 1520 0 sw_n2
rlabel metal2 12190 1520 12190 1520 0 sw_n3
rlabel metal2 10902 823 10902 823 0 sw_n4
rlabel metal1 9706 3366 9706 3366 0 sw_n5
rlabel metal1 4738 2822 4738 2822 0 sw_n6
rlabel metal2 3174 1520 3174 1520 0 sw_n7
rlabel metal2 1886 1520 1886 1520 0 sw_n8
rlabel metal2 21206 1520 21206 1520 0 sw_n_sp1
rlabel metal2 19918 1520 19918 1520 0 sw_n_sp2
rlabel metal2 16054 1520 16054 1520 0 sw_n_sp3
rlabel metal2 14766 1520 14766 1520 0 sw_n_sp4
rlabel metal2 13478 1520 13478 1520 0 sw_n_sp5
rlabel metal2 8326 1520 8326 1520 0 sw_n_sp6
rlabel metal2 7038 1520 7038 1520 0 sw_n_sp7
rlabel metal2 5750 1520 5750 1520 0 sw_n_sp8
rlabel metal2 598 1520 598 1520 0 sw_n_sp9
rlabel metal1 19044 21658 19044 21658 0 sw_p1
rlabel metal2 17618 22491 17618 22491 0 sw_p2
rlabel metal1 12236 21590 12236 21590 0 sw_p3
rlabel metal2 10757 23324 10757 23324 0 sw_p4
rlabel metal1 9660 21590 9660 21590 0 sw_p5
rlabel metal2 4515 23324 4515 23324 0 sw_p6
rlabel metal1 3588 21658 3588 21658 0 sw_p7
rlabel metal2 1978 22457 1978 22457 0 sw_p8
rlabel metal1 20700 21114 20700 21114 0 sw_p_sp1
rlabel metal2 20102 22491 20102 22491 0 sw_p_sp2
rlabel metal2 16054 22484 16054 22484 0 sw_p_sp3
rlabel metal1 14996 21658 14996 21658 0 sw_p_sp4
rlabel metal1 13892 21658 13892 21658 0 sw_p_sp5
rlabel metal1 8740 21658 8740 21658 0 sw_p_sp6
rlabel metal1 7176 21658 7176 21658 0 sw_p_sp7
rlabel metal1 6164 21658 6164 21658 0 sw_p_sp8
rlabel metal1 1104 21658 1104 21658 0 sw_p_sp9
rlabel metal1 1426 21114 1426 21114 0 sw_sample
rlabel metal2 17986 19856 17986 19856 0 x1/cycle0
rlabel metal1 16606 15606 16606 15606 0 x1/cycle1
rlabel metal1 10672 6630 10672 6630 0 x1/cycle10
rlabel metal1 3082 19414 3082 19414 0 x1/cycle11
rlabel metal1 15870 5780 15870 5780 0 x1/cycle12
rlabel metal1 16192 5270 16192 5270 0 x1/cycle13
rlabel metal2 17342 7820 17342 7820 0 x1/cycle14
rlabel metal1 17434 7276 17434 7276 0 x1/cycle15
rlabel metal1 14306 17170 14306 17170 0 x1/cycle2
rlabel metal1 14030 14450 14030 14450 0 x1/cycle3
rlabel metal1 16629 12818 16629 12818 0 x1/cycle4
rlabel metal2 12374 10370 12374 10370 0 x1/cycle5
rlabel metal1 14398 10200 14398 10200 0 x1/cycle6
rlabel metal1 4554 2482 4554 2482 0 x1/cycle7
rlabel metal1 8602 5780 8602 5780 0 x1/cycle8
rlabel metal2 3818 4794 3818 4794 0 x1/cycle9
rlabel metal2 17710 7956 17710 7956 0 x1/net1
rlabel metal1 18124 8466 18124 8466 0 x1/net2
rlabel metal1 18354 7854 18354 7854 0 x1/net3
rlabel metal2 18630 7582 18630 7582 0 x1/net4
rlabel metal1 1794 13294 1794 13294 0 x1/net5
rlabel metal2 2254 13634 2254 13634 0 x1/net6
rlabel metal2 17710 14688 17710 14688 0 x1/raw_bit1
rlabel metal2 12282 4998 12282 4998 0 x1/raw_bit10
rlabel metal1 13524 5542 13524 5542 0 x1/raw_bit11
rlabel metal1 14490 3162 14490 3162 0 x1/raw_bit12
rlabel metal1 18814 4046 18814 4046 0 x1/raw_bit13
rlabel metal1 18453 14994 18453 14994 0 x1/raw_bit2
rlabel metal1 16790 15606 16790 15606 0 x1/raw_bit3
rlabel metal2 17434 10336 17434 10336 0 x1/raw_bit4
rlabel metal2 18446 12410 18446 12410 0 x1/raw_bit5
rlabel metal2 17158 10914 17158 10914 0 x1/raw_bit6
rlabel metal1 16514 10064 16514 10064 0 x1/raw_bit7
rlabel metal2 14398 5372 14398 5372 0 x1/raw_bit8
rlabel metal1 14306 5787 14306 5787 0 x1/raw_bit9
rlabel metal1 17986 6290 17986 6290 0 x1/raw_bit_clr
rlabel metal1 15042 9928 15042 9928 0 x1/vcmp_buf
rlabel metal1 17572 15130 17572 15130 0 x1/x1/net1
rlabel metal1 18722 8534 18722 8534 0 x1/x1/net10
rlabel metal1 17434 5576 17434 5576 0 x1/x1/net11
rlabel metal2 18906 6052 18906 6052 0 x1/x1/net12
rlabel metal1 14076 5338 14076 5338 0 x1/x1/net13
rlabel metal1 16767 5270 16767 5270 0 x1/x1/net14
rlabel metal2 14122 4930 14122 4930 0 x1/x1/net15
rlabel metal2 18814 4964 18814 4964 0 x1/x1/net16
rlabel metal1 18722 15062 18722 15062 0 x1/x1/net2
rlabel metal2 17066 14722 17066 14722 0 x1/x1/net3
rlabel metal1 18676 13974 18676 13974 0 x1/x1/net4
rlabel metal2 18906 11934 18906 11934 0 x1/x1/net5
rlabel metal2 17250 13464 17250 13464 0 x1/x1/net6
rlabel metal1 17388 10778 17388 10778 0 x1/x1/net7
rlabel metal1 18722 10710 18722 10710 0 x1/x1/net8
rlabel metal1 17204 10234 17204 10234 0 x1/x1/net9
rlabel metal1 18699 20502 18699 20502 0 x1/x2/net1
rlabel metal2 16054 18564 16054 18564 0 x1/x2/net10
rlabel metal1 17112 3026 17112 3026 0 x1/x2/net11
rlabel metal1 15410 3570 15410 3570 0 x1/x2/net12
rlabel metal1 14352 14314 14352 14314 0 x1/x2/net13
rlabel metal2 15410 13770 15410 13770 0 x1/x2/net14
rlabel metal1 13685 13838 13685 13838 0 x1/x2/net15
rlabel metal2 13294 15232 13294 15232 0 x1/x2/net16
rlabel metal2 14030 13430 14030 13430 0 x1/x2/net17
rlabel metal1 14053 10778 14053 10778 0 x1/x2/net18
rlabel metal1 11707 15402 11707 15402 0 x1/x2/net19
rlabel metal2 19642 19176 19642 19176 0 x1/x2/net2
rlabel metal1 10925 20978 10925 20978 0 x1/x2/net20
rlabel metal2 13110 13702 13110 13702 0 x1/x2/net21
rlabel metal2 14490 10438 14490 10438 0 x1/x2/net22
rlabel metal1 11477 11322 11477 11322 0 x1/x2/net23
rlabel metal2 12466 13770 12466 13770 0 x1/x2/net24
rlabel metal2 9614 20604 9614 20604 0 x1/x2/net25
rlabel metal1 8533 17170 8533 17170 0 x1/x2/net26
rlabel metal1 13202 10098 13202 10098 0 x1/x2/net27
rlabel metal1 8970 17102 8970 17102 0 x1/x2/net28
rlabel metal1 11086 10778 11086 10778 0 x1/x2/net29
rlabel metal1 18837 17646 18837 17646 0 x1/x2/net3
rlabel metal1 11408 13498 11408 13498 0 x1/x2/net30
rlabel metal1 6923 6426 6923 6426 0 x1/x2/net31
rlabel metal1 7820 3706 7820 3706 0 x1/x2/net32
rlabel metal2 8234 3740 8234 3740 0 x1/x2/net33
rlabel metal2 4738 9758 4738 9758 0 x1/x2/net34
rlabel metal1 5658 5338 5658 5338 0 x1/x2/net35
rlabel metal1 5267 4794 5267 4794 0 x1/x2/net36
rlabel metal1 4370 9010 4370 9010 0 x1/x2/net37
rlabel metal1 3496 14994 3496 14994 0 x1/x2/net38
rlabel metal1 8430 4114 8430 4114 0 x1/x2/net39
rlabel metal2 18262 19550 18262 19550 0 x1/x2/net4
rlabel metal1 5302 4590 5302 4590 0 x1/x2/net40
rlabel metal1 5175 7854 5175 7854 0 x1/x2/net41
rlabel metal1 4784 7718 4784 7718 0 x1/x2/net42
rlabel via1 1909 17306 1909 17306 0 x1/x2/net43
rlabel metal1 1863 15130 1863 15130 0 x1/x2/net44
rlabel metal2 1426 5372 1426 5372 0 x1/x2/net45
rlabel metal1 2346 15538 2346 15538 0 x1/x2/net46
rlabel metal1 5364 7854 5364 7854 0 x1/x2/net47
rlabel metal1 2990 2958 2990 2958 0 x1/x2/net48
rlabel metal2 2898 19108 2898 19108 0 x1/x2/net49
rlabel metal2 18814 18870 18814 18870 0 x1/x2/net5
rlabel metal2 17158 16898 17158 16898 0 x1/x2/net50
rlabel metal1 16675 17170 16675 17170 0 x1/x2/net51
rlabel metal1 17204 17170 17204 17170 0 x1/x2/net52
rlabel metal2 15686 16796 15686 16796 0 x1/x2/net53
rlabel metal2 15686 18224 15686 18224 0 x1/x2/net54
rlabel metal1 14122 17306 14122 17306 0 x1/x2/net55
rlabel metal1 15410 18190 15410 18190 0 x1/x2/net56
rlabel metal1 14168 17714 14168 17714 0 x1/x2/net57
rlabel via1 12177 12818 12177 12818 0 x1/x2/net58
rlabel metal1 11592 12818 11592 12818 0 x1/x2/net59
rlabel metal1 17043 18734 17043 18734 0 x1/x2/net6
rlabel metal1 12926 13260 12926 13260 0 x1/x2/net60
rlabel metal2 10626 12988 10626 12988 0 x1/x2/net61
rlabel metal1 13524 10166 13524 10166 0 x1/x2/net62
rlabel metal1 13202 9418 13202 9418 0 x1/x2/net63
rlabel metal1 14122 10166 14122 10166 0 x1/x2/net64
rlabel metal1 11546 10098 11546 10098 0 x1/x2/net65
rlabel metal2 10534 10234 10534 10234 0 x1/x2/net66
rlabel metal1 8970 10778 8970 10778 0 x1/x2/net67
rlabel metal2 9798 10846 9798 10846 0 x1/x2/net68
rlabel metal2 9154 10404 9154 10404 0 x1/x2/net69
rlabel metal1 17181 20978 17181 20978 0 x1/x2/net7
rlabel metal1 8400 4590 8400 4590 0 x1/x2/net70
rlabel metal1 7314 4590 7314 4590 0 x1/x2/net71
rlabel metal1 7820 4590 7820 4590 0 x1/x2/net72
rlabel metal1 6394 5066 6394 5066 0 x1/x2/net73
rlabel metal1 5152 5338 5152 5338 0 x1/x2/net74
rlabel metal1 4140 4590 4140 4590 0 x1/x2/net75
rlabel metal2 4462 5236 4462 5236 0 x1/x2/net76
rlabel metal1 3404 5270 3404 5270 0 x1/x2/net77
rlabel metal1 4232 7922 4232 7922 0 x1/x2/net78
rlabel metal1 2530 7752 2530 7752 0 x1/x2/net79
rlabel metal1 15709 19890 15709 19890 0 x1/x2/net8
rlabel metal1 3450 7820 3450 7820 0 x1/x2/net80
rlabel metal1 3036 6970 3036 6970 0 x1/x2/net81
rlabel metal2 18078 17476 18078 17476 0 x1/x2/net9
rlabel metal2 12558 13124 12558 13124 0 x1/x2/x119/net1
rlabel metal1 17457 16762 17457 16762 0 x1/x2/x16/net1
rlabel metal1 15157 18190 15157 18190 0 x1/x2/x17/net1
rlabel metal1 13455 9690 13455 9690 0 x1/x2/x35/net1
rlabel via1 9913 10234 9913 10234 0 x1/x2/x36/net1
rlabel metal1 8211 4590 8211 4590 0 x1/x2/x39/net1
rlabel metal1 4991 5678 4991 5678 0 x1/x2/x62/net1
rlabel metal1 3749 7854 3749 7854 0 x1/x2/x63/net1
rlabel metal1 9660 18326 9660 18326 0 x1/x3/count_net
rlabel via1 8993 20026 8993 20026 0 x1/x3/johnson_counter_loop
rlabel metal1 4508 20366 4508 20366 0 x1/x3/net1
rlabel metal1 12880 19482 12880 19482 0 x1/x3/net10
rlabel metal2 13938 20196 13938 20196 0 x1/x3/net11
rlabel metal1 14628 20570 14628 20570 0 x1/x3/net12
rlabel metal2 15226 20332 15226 20332 0 x1/x3/net13
rlabel metal1 7176 20026 7176 20026 0 x1/x3/net14
rlabel metal1 4462 20026 4462 20026 0 x1/x3/net15
rlabel metal1 4554 20910 4554 20910 0 x1/x3/net16
rlabel via1 9136 19822 9136 19822 0 x1/x3/net17
rlabel metal2 3542 17340 3542 17340 0 x1/x3/net18
rlabel metal1 3312 16626 3312 16626 0 x1/x3/net19
rlabel metal1 5198 19414 5198 19414 0 x1/x3/net2
rlabel metal2 3174 16762 3174 16762 0 x1/x3/net20
rlabel metal1 2944 16626 2944 16626 0 x1/x3/net21
rlabel metal2 2438 10812 2438 10812 0 x1/x3/net22
rlabel metal2 2346 10234 2346 10234 0 x1/x3/net23
rlabel metal2 2990 9758 2990 9758 0 x1/x3/net24
rlabel metal2 4370 18904 4370 18904 0 x1/x3/net3
rlabel metal1 5796 18394 5796 18394 0 x1/x3/net4
rlabel metal1 6670 17714 6670 17714 0 x1/x3/net5
rlabel metal2 7866 18020 7866 18020 0 x1/x3/net6
rlabel metal1 8832 18394 8832 18394 0 x1/x3/net7
rlabel metal1 10856 18394 10856 18394 0 x1/x3/net8
rlabel metal1 11960 18938 11960 18938 0 x1/x3/net9
rlabel metal2 8050 15844 8050 15844 0 x1/x4/net1
rlabel metal1 9476 7446 9476 7446 0 x1/x4/net10
rlabel metal1 10672 7514 10672 7514 0 x1/x4/net11
rlabel metal2 11914 8262 11914 8262 0 x1/x4/net12
rlabel metal1 14168 6766 14168 6766 0 x1/x4/net13
rlabel metal1 14858 7514 14858 7514 0 x1/x4/net14
rlabel metal2 16606 7650 16606 7650 0 x1/x4/net15
rlabel metal2 5198 14756 5198 14756 0 x1/x4/net16
rlabel metal2 6394 15436 6394 15436 0 x1/x4/net17
rlabel metal1 6946 16014 6946 16014 0 x1/x4/net18
rlabel metal1 6072 16082 6072 16082 0 x1/x4/net19
rlabel metal1 9706 16048 9706 16048 0 x1/x4/net2
rlabel metal1 9430 14892 9430 14892 0 x1/x4/net20
rlabel metal1 8786 15538 8786 15538 0 x1/x4/net21
rlabel metal2 8418 15300 8418 15300 0 x1/x4/net22
rlabel metal1 8096 14994 8096 14994 0 x1/x4/net23
rlabel metal2 16330 8126 16330 8126 0 x1/x4/net24
rlabel metal1 14398 7922 14398 7922 0 x1/x4/net25
rlabel metal1 13202 7276 13202 7276 0 x1/x4/net26
rlabel metal2 12006 8092 12006 8092 0 x1/x4/net27
rlabel metal1 10028 7922 10028 7922 0 x1/x4/net28
rlabel metal2 9154 7548 9154 7548 0 x1/x4/net29
rlabel metal1 10350 15334 10350 15334 0 x1/x4/net3
rlabel metal1 7774 8364 7774 8364 0 x1/x4/net30
rlabel metal1 6624 7922 6624 7922 0 x1/x4/net31
rlabel metal2 6394 10812 6394 10812 0 x1/x4/net32
rlabel metal2 6210 11356 6210 11356 0 x1/x4/net33
rlabel metal1 8234 12716 8234 12716 0 x1/x4/net34
rlabel metal2 7866 13668 7866 13668 0 x1/x4/net35
rlabel metal1 7636 13294 7636 13294 0 x1/x4/net36
rlabel metal1 6118 11730 6118 11730 0 x1/x4/net37
rlabel metal1 7268 7514 7268 7514 0 x1/x4/net38
rlabel metal1 9200 7990 9200 7990 0 x1/x4/net39
rlabel metal2 11178 14280 11178 14280 0 x1/x4/net4
rlabel metal2 12466 7990 12466 7990 0 x1/x4/net40
rlabel metal1 13754 8466 13754 8466 0 x1/x4/net41
rlabel metal2 12558 7888 12558 7888 0 x1/x4/net42
rlabel metal1 8924 16762 8924 16762 0 x1/x4/net43
rlabel metal2 9890 16388 9890 16388 0 x1/x4/net44
rlabel metal2 11270 15878 11270 15878 0 x1/x4/net45
rlabel metal1 11730 15096 11730 15096 0 x1/x4/net46
rlabel metal1 9752 13294 9752 13294 0 x1/x4/net47
rlabel metal1 11362 11152 11362 11152 0 x1/x4/net48
rlabel metal2 7958 10438 7958 10438 0 x1/x4/net49
rlabel metal1 9016 13294 9016 13294 0 x1/x4/net5
rlabel metal1 7084 8874 7084 8874 0 x1/x4/net50
rlabel metal2 8786 6154 8786 6154 0 x1/x4/net51
rlabel metal2 9614 5644 9614 5644 0 x1/x4/net52
rlabel metal2 10994 6970 10994 6970 0 x1/x4/net53
rlabel metal2 11822 7854 11822 7854 0 x1/x4/net54
rlabel metal1 15088 6630 15088 6630 0 x1/x4/net55
rlabel metal2 15502 7990 15502 7990 0 x1/x4/net56
rlabel metal1 17066 7514 17066 7514 0 x1/x4/net57
rlabel metal2 17986 7854 17986 7854 0 x1/x4/net58
rlabel metal1 18308 8058 18308 8058 0 x1/x4/net59
rlabel metal1 9936 12614 9936 12614 0 x1/x4/net6
rlabel metal1 4531 16558 4531 16558 0 x1/x4/net60
rlabel metal2 5014 15946 5014 15946 0 x1/x4/net61
rlabel metal1 7820 10030 7820 10030 0 x1/x4/net7
rlabel metal1 7866 8942 7866 8942 0 x1/x4/net8
rlabel metal1 8556 8058 8556 8058 0 x1/x4/net9
rlabel metal1 7360 15470 7360 15470 0 x1/x4/reset_b
rlabel metal1 2898 11628 2898 11628 0 x2/net1
rlabel metal1 4692 12206 4692 12206 0 x2/net10
rlabel metal1 5336 13294 5336 13294 0 x2/net11
rlabel metal1 2576 11730 2576 11730 0 x2/net2
rlabel metal1 2622 11832 2622 11832 0 x2/net3
rlabel metal1 3358 11730 3358 11730 0 x2/net4
rlabel metal1 3864 11730 3864 11730 0 x2/net5
rlabel metal1 4600 11866 4600 11866 0 x2/net6
rlabel metal2 4922 13124 4922 13124 0 x2/net7
rlabel metal1 4876 12818 4876 12818 0 x2/net8
rlabel metal1 4968 12410 4968 12410 0 x2/net9
<< properties >>
string FIXED_BBOX 0 0 21880 24024
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1754794521
<< error_p >>
rect -653 163 -595 169
rect -461 163 -403 169
rect -269 163 -211 169
rect -77 163 -19 169
rect 115 163 173 169
rect 307 163 365 169
rect 499 163 557 169
rect 691 163 749 169
rect -653 129 -641 163
rect -461 129 -449 163
rect -269 129 -257 163
rect -77 129 -65 163
rect 115 129 127 163
rect 307 129 319 163
rect 499 129 511 163
rect 691 129 703 163
rect -653 123 -595 129
rect -461 123 -403 129
rect -269 123 -211 129
rect -77 123 -19 129
rect 115 123 173 129
rect 307 123 365 129
rect 499 123 557 129
rect 691 123 749 129
rect -791 62 -745 74
rect -599 62 -553 74
rect -407 62 -361 74
rect -215 62 -169 74
rect -23 62 23 74
rect 169 62 215 74
rect 361 62 407 74
rect 553 62 599 74
rect 745 62 791 74
rect -791 15 -785 62
rect -599 15 -593 62
rect -407 15 -401 62
rect -215 15 -209 62
rect -23 15 -17 62
rect 169 15 175 62
rect 361 15 367 62
rect 553 15 559 62
rect 745 15 751 62
rect -791 3 -745 15
rect -599 3 -553 15
rect -407 3 -361 15
rect -215 3 -169 15
rect -23 3 23 15
rect 169 3 215 15
rect 361 3 407 15
rect 553 3 599 15
rect 745 3 791 15
rect -695 -15 -649 -3
rect -503 -15 -457 -3
rect -311 -15 -265 -3
rect -119 -15 -73 -3
rect 73 -15 119 -3
rect 265 -15 311 -3
rect 457 -15 503 -3
rect 649 -15 695 -3
rect -695 -62 -689 -15
rect -503 -62 -497 -15
rect -311 -62 -305 -15
rect -119 -62 -113 -15
rect 73 -62 79 -15
rect 265 -62 271 -15
rect 457 -62 463 -15
rect 649 -62 655 -15
rect -695 -74 -649 -62
rect -503 -74 -457 -62
rect -311 -74 -265 -62
rect -119 -74 -73 -62
rect 73 -74 119 -62
rect 265 -74 311 -62
rect 457 -74 503 -62
rect 649 -74 695 -62
rect -749 -129 -691 -123
rect -557 -129 -499 -123
rect -365 -129 -307 -123
rect -173 -129 -115 -123
rect 19 -129 77 -123
rect 211 -129 269 -123
rect 403 -129 461 -123
rect 595 -129 653 -123
rect -749 -163 -737 -129
rect -557 -163 -545 -129
rect -365 -163 -353 -129
rect -173 -163 -161 -129
rect 19 -163 31 -129
rect 211 -163 223 -129
rect 403 -163 415 -129
rect 595 -163 607 -129
rect -749 -169 -691 -163
rect -557 -169 -499 -163
rect -365 -169 -307 -163
rect -173 -169 -115 -163
rect 19 -169 77 -163
rect 211 -169 269 -163
rect 403 -169 461 -163
rect 595 -169 653 -163
<< nmos >>
rect -735 -91 -705 91
rect -639 -91 -609 91
rect -543 -91 -513 91
rect -447 -91 -417 91
rect -351 -91 -321 91
rect -255 -91 -225 91
rect -159 -91 -129 91
rect -63 -91 -33 91
rect 33 -91 63 91
rect 129 -91 159 91
rect 225 -91 255 91
rect 321 -91 351 91
rect 417 -91 447 91
rect 513 -91 543 91
rect 609 -91 639 91
rect 705 -91 735 91
<< ndiff >>
rect -797 79 -735 91
rect -797 -79 -785 79
rect -751 -79 -735 79
rect -797 -91 -735 -79
rect -705 79 -639 91
rect -705 -79 -689 79
rect -655 -79 -639 79
rect -705 -91 -639 -79
rect -609 79 -543 91
rect -609 -79 -593 79
rect -559 -79 -543 79
rect -609 -91 -543 -79
rect -513 79 -447 91
rect -513 -79 -497 79
rect -463 -79 -447 79
rect -513 -91 -447 -79
rect -417 79 -351 91
rect -417 -79 -401 79
rect -367 -79 -351 79
rect -417 -91 -351 -79
rect -321 79 -255 91
rect -321 -79 -305 79
rect -271 -79 -255 79
rect -321 -91 -255 -79
rect -225 79 -159 91
rect -225 -79 -209 79
rect -175 -79 -159 79
rect -225 -91 -159 -79
rect -129 79 -63 91
rect -129 -79 -113 79
rect -79 -79 -63 79
rect -129 -91 -63 -79
rect -33 79 33 91
rect -33 -79 -17 79
rect 17 -79 33 79
rect -33 -91 33 -79
rect 63 79 129 91
rect 63 -79 79 79
rect 113 -79 129 79
rect 63 -91 129 -79
rect 159 79 225 91
rect 159 -79 175 79
rect 209 -79 225 79
rect 159 -91 225 -79
rect 255 79 321 91
rect 255 -79 271 79
rect 305 -79 321 79
rect 255 -91 321 -79
rect 351 79 417 91
rect 351 -79 367 79
rect 401 -79 417 79
rect 351 -91 417 -79
rect 447 79 513 91
rect 447 -79 463 79
rect 497 -79 513 79
rect 447 -91 513 -79
rect 543 79 609 91
rect 543 -79 559 79
rect 593 -79 609 79
rect 543 -91 609 -79
rect 639 79 705 91
rect 639 -79 655 79
rect 689 -79 705 79
rect 639 -91 705 -79
rect 735 79 797 91
rect 735 -79 751 79
rect 785 -79 797 79
rect 735 -91 797 -79
<< ndiffc >>
rect -785 -79 -751 79
rect -689 -79 -655 79
rect -593 -79 -559 79
rect -497 -79 -463 79
rect -401 -79 -367 79
rect -305 -79 -271 79
rect -209 -79 -175 79
rect -113 -79 -79 79
rect -17 -79 17 79
rect 79 -79 113 79
rect 175 -79 209 79
rect 271 -79 305 79
rect 367 -79 401 79
rect 463 -79 497 79
rect 559 -79 593 79
rect 655 -79 689 79
rect 751 -79 785 79
<< poly >>
rect -657 163 -591 179
rect -657 129 -641 163
rect -607 129 -591 163
rect -735 91 -705 117
rect -657 113 -591 129
rect -465 163 -399 179
rect -465 129 -449 163
rect -415 129 -399 163
rect -639 91 -609 113
rect -543 91 -513 117
rect -465 113 -399 129
rect -273 163 -207 179
rect -273 129 -257 163
rect -223 129 -207 163
rect -447 91 -417 113
rect -351 91 -321 117
rect -273 113 -207 129
rect -81 163 -15 179
rect -81 129 -65 163
rect -31 129 -15 163
rect -255 91 -225 113
rect -159 91 -129 117
rect -81 113 -15 129
rect 111 163 177 179
rect 111 129 127 163
rect 161 129 177 163
rect -63 91 -33 113
rect 33 91 63 117
rect 111 113 177 129
rect 303 163 369 179
rect 303 129 319 163
rect 353 129 369 163
rect 129 91 159 113
rect 225 91 255 117
rect 303 113 369 129
rect 495 163 561 179
rect 495 129 511 163
rect 545 129 561 163
rect 321 91 351 113
rect 417 91 447 117
rect 495 113 561 129
rect 687 163 753 179
rect 687 129 703 163
rect 737 129 753 163
rect 513 91 543 113
rect 609 91 639 117
rect 687 113 753 129
rect 705 91 735 113
rect -735 -113 -705 -91
rect -753 -129 -687 -113
rect -639 -117 -609 -91
rect -543 -113 -513 -91
rect -753 -163 -737 -129
rect -703 -163 -687 -129
rect -753 -179 -687 -163
rect -561 -129 -495 -113
rect -447 -117 -417 -91
rect -351 -113 -321 -91
rect -561 -163 -545 -129
rect -511 -163 -495 -129
rect -561 -179 -495 -163
rect -369 -129 -303 -113
rect -255 -117 -225 -91
rect -159 -113 -129 -91
rect -369 -163 -353 -129
rect -319 -163 -303 -129
rect -369 -179 -303 -163
rect -177 -129 -111 -113
rect -63 -117 -33 -91
rect 33 -113 63 -91
rect -177 -163 -161 -129
rect -127 -163 -111 -129
rect -177 -179 -111 -163
rect 15 -129 81 -113
rect 129 -117 159 -91
rect 225 -113 255 -91
rect 15 -163 31 -129
rect 65 -163 81 -129
rect 15 -179 81 -163
rect 207 -129 273 -113
rect 321 -117 351 -91
rect 417 -113 447 -91
rect 207 -163 223 -129
rect 257 -163 273 -129
rect 207 -179 273 -163
rect 399 -129 465 -113
rect 513 -117 543 -91
rect 609 -113 639 -91
rect 399 -163 415 -129
rect 449 -163 465 -129
rect 399 -179 465 -163
rect 591 -129 657 -113
rect 705 -117 735 -91
rect 591 -163 607 -129
rect 641 -163 657 -129
rect 591 -179 657 -163
<< polycont >>
rect -641 129 -607 163
rect -449 129 -415 163
rect -257 129 -223 163
rect -65 129 -31 163
rect 127 129 161 163
rect 319 129 353 163
rect 511 129 545 163
rect 703 129 737 163
rect -737 -163 -703 -129
rect -545 -163 -511 -129
rect -353 -163 -319 -129
rect -161 -163 -127 -129
rect 31 -163 65 -129
rect 223 -163 257 -129
rect 415 -163 449 -129
rect 607 -163 641 -129
<< locali >>
rect -657 129 -641 163
rect -607 129 -591 163
rect -465 129 -449 163
rect -415 129 -399 163
rect -273 129 -257 163
rect -223 129 -207 163
rect -81 129 -65 163
rect -31 129 -15 163
rect 111 129 127 163
rect 161 129 177 163
rect 303 129 319 163
rect 353 129 369 163
rect 495 129 511 163
rect 545 129 561 163
rect 687 129 703 163
rect 737 129 753 163
rect -785 79 -751 95
rect -785 -95 -751 -79
rect -689 79 -655 95
rect -689 -95 -655 -79
rect -593 79 -559 95
rect -593 -95 -559 -79
rect -497 79 -463 95
rect -497 -95 -463 -79
rect -401 79 -367 95
rect -401 -95 -367 -79
rect -305 79 -271 95
rect -305 -95 -271 -79
rect -209 79 -175 95
rect -209 -95 -175 -79
rect -113 79 -79 95
rect -113 -95 -79 -79
rect -17 79 17 95
rect -17 -95 17 -79
rect 79 79 113 95
rect 79 -95 113 -79
rect 175 79 209 95
rect 175 -95 209 -79
rect 271 79 305 95
rect 271 -95 305 -79
rect 367 79 401 95
rect 367 -95 401 -79
rect 463 79 497 95
rect 463 -95 497 -79
rect 559 79 593 95
rect 559 -95 593 -79
rect 655 79 689 95
rect 655 -95 689 -79
rect 751 79 785 95
rect 751 -95 785 -79
rect -753 -163 -737 -129
rect -703 -163 -687 -129
rect -561 -163 -545 -129
rect -511 -163 -495 -129
rect -369 -163 -353 -129
rect -319 -163 -303 -129
rect -177 -163 -161 -129
rect -127 -163 -111 -129
rect 15 -163 31 -129
rect 65 -163 81 -129
rect 207 -163 223 -129
rect 257 -163 273 -129
rect 399 -163 415 -129
rect 449 -163 465 -129
rect 591 -163 607 -129
rect 641 -163 657 -129
<< viali >>
rect -641 129 -607 163
rect -449 129 -415 163
rect -257 129 -223 163
rect -65 129 -31 163
rect 127 129 161 163
rect 319 129 353 163
rect 511 129 545 163
rect 703 129 737 163
rect -785 15 -751 62
rect -689 -62 -655 -15
rect -593 15 -559 62
rect -497 -62 -463 -15
rect -401 15 -367 62
rect -305 -62 -271 -15
rect -209 15 -175 62
rect -113 -62 -79 -15
rect -17 15 17 62
rect 79 -62 113 -15
rect 175 15 209 62
rect 271 -62 305 -15
rect 367 15 401 62
rect 463 -62 497 -15
rect 559 15 593 62
rect 655 -62 689 -15
rect 751 15 785 62
rect -737 -163 -703 -129
rect -545 -163 -511 -129
rect -353 -163 -319 -129
rect -161 -163 -127 -129
rect 31 -163 65 -129
rect 223 -163 257 -129
rect 415 -163 449 -129
rect 607 -163 641 -129
<< metal1 >>
rect -653 163 -595 169
rect -653 129 -641 163
rect -607 129 -595 163
rect -653 123 -595 129
rect -461 163 -403 169
rect -461 129 -449 163
rect -415 129 -403 163
rect -461 123 -403 129
rect -269 163 -211 169
rect -269 129 -257 163
rect -223 129 -211 163
rect -269 123 -211 129
rect -77 163 -19 169
rect -77 129 -65 163
rect -31 129 -19 163
rect -77 123 -19 129
rect 115 163 173 169
rect 115 129 127 163
rect 161 129 173 163
rect 115 123 173 129
rect 307 163 365 169
rect 307 129 319 163
rect 353 129 365 163
rect 307 123 365 129
rect 499 163 557 169
rect 499 129 511 163
rect 545 129 557 163
rect 499 123 557 129
rect 691 163 749 169
rect 691 129 703 163
rect 737 129 749 163
rect 691 123 749 129
rect -791 62 -745 74
rect -791 15 -785 62
rect -751 15 -745 62
rect -791 3 -745 15
rect -599 62 -553 74
rect -599 15 -593 62
rect -559 15 -553 62
rect -599 3 -553 15
rect -407 62 -361 74
rect -407 15 -401 62
rect -367 15 -361 62
rect -407 3 -361 15
rect -215 62 -169 74
rect -215 15 -209 62
rect -175 15 -169 62
rect -215 3 -169 15
rect -23 62 23 74
rect -23 15 -17 62
rect 17 15 23 62
rect -23 3 23 15
rect 169 62 215 74
rect 169 15 175 62
rect 209 15 215 62
rect 169 3 215 15
rect 361 62 407 74
rect 361 15 367 62
rect 401 15 407 62
rect 361 3 407 15
rect 553 62 599 74
rect 553 15 559 62
rect 593 15 599 62
rect 553 3 599 15
rect 745 62 791 74
rect 745 15 751 62
rect 785 15 791 62
rect 745 3 791 15
rect -695 -15 -649 -3
rect -695 -62 -689 -15
rect -655 -62 -649 -15
rect -695 -74 -649 -62
rect -503 -15 -457 -3
rect -503 -62 -497 -15
rect -463 -62 -457 -15
rect -503 -74 -457 -62
rect -311 -15 -265 -3
rect -311 -62 -305 -15
rect -271 -62 -265 -15
rect -311 -74 -265 -62
rect -119 -15 -73 -3
rect -119 -62 -113 -15
rect -79 -62 -73 -15
rect -119 -74 -73 -62
rect 73 -15 119 -3
rect 73 -62 79 -15
rect 113 -62 119 -15
rect 73 -74 119 -62
rect 265 -15 311 -3
rect 265 -62 271 -15
rect 305 -62 311 -15
rect 265 -74 311 -62
rect 457 -15 503 -3
rect 457 -62 463 -15
rect 497 -62 503 -15
rect 457 -74 503 -62
rect 649 -15 695 -3
rect 649 -62 655 -15
rect 689 -62 695 -15
rect 649 -74 695 -62
rect -749 -129 -691 -123
rect -749 -163 -737 -129
rect -703 -163 -691 -129
rect -749 -169 -691 -163
rect -557 -129 -499 -123
rect -557 -163 -545 -129
rect -511 -163 -499 -129
rect -557 -169 -499 -163
rect -365 -129 -307 -123
rect -365 -163 -353 -129
rect -319 -163 -307 -129
rect -365 -169 -307 -163
rect -173 -129 -115 -123
rect -173 -163 -161 -129
rect -127 -163 -115 -129
rect -173 -169 -115 -163
rect 19 -129 77 -123
rect 19 -163 31 -129
rect 65 -163 77 -129
rect 19 -169 77 -163
rect 211 -129 269 -123
rect 211 -163 223 -129
rect 257 -163 269 -129
rect 211 -169 269 -163
rect 403 -129 461 -123
rect 403 -163 415 -129
rect 449 -163 461 -129
rect 403 -169 461 -163
rect 595 -129 653 -123
rect 595 -163 607 -129
rect 641 -163 653 -129
rect 595 -169 653 -163
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.91 l 0.15 m 1 nf 16 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc +30 viadrn -30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

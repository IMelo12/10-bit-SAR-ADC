** sch_path: /home/ttuser/Documents/SARADC/xschem/cap16/cap16.sch
**.subckt cap16 bottom top
*.ipin bottom
*.ipin top
XC12 top bottom sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=16 m=16
**.ends
.end

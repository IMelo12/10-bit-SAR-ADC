magic
tech sky130A
magscale 1 2
timestamp 1754899980
<< metal3 >>
rect -1492 10412 -120 10440
rect -1492 9388 -204 10412
rect -140 9388 -120 10412
rect -1492 9360 -120 9388
rect 120 10412 1492 10440
rect 120 9388 1408 10412
rect 1472 9388 1492 10412
rect 120 9360 1492 9388
rect -1492 9092 -120 9120
rect -1492 8068 -204 9092
rect -140 8068 -120 9092
rect -1492 8040 -120 8068
rect 120 9092 1492 9120
rect 120 8068 1408 9092
rect 1472 8068 1492 9092
rect 120 8040 1492 8068
rect -1492 7772 -120 7800
rect -1492 6748 -204 7772
rect -140 6748 -120 7772
rect -1492 6720 -120 6748
rect 120 7772 1492 7800
rect 120 6748 1408 7772
rect 1472 6748 1492 7772
rect 120 6720 1492 6748
rect -1492 6452 -120 6480
rect -1492 5428 -204 6452
rect -140 5428 -120 6452
rect -1492 5400 -120 5428
rect 120 6452 1492 6480
rect 120 5428 1408 6452
rect 1472 5428 1492 6452
rect 120 5400 1492 5428
rect -1492 5132 -120 5160
rect -1492 4108 -204 5132
rect -140 4108 -120 5132
rect -1492 4080 -120 4108
rect 120 5132 1492 5160
rect 120 4108 1408 5132
rect 1472 4108 1492 5132
rect 120 4080 1492 4108
rect -1492 3812 -120 3840
rect -1492 2788 -204 3812
rect -140 2788 -120 3812
rect -1492 2760 -120 2788
rect 120 3812 1492 3840
rect 120 2788 1408 3812
rect 1472 2788 1492 3812
rect 120 2760 1492 2788
rect -1492 2492 -120 2520
rect -1492 1468 -204 2492
rect -140 1468 -120 2492
rect -1492 1440 -120 1468
rect 120 2492 1492 2520
rect 120 1468 1408 2492
rect 1472 1468 1492 2492
rect 120 1440 1492 1468
rect -1492 1172 -120 1200
rect -1492 148 -204 1172
rect -140 148 -120 1172
rect -1492 120 -120 148
rect 120 1172 1492 1200
rect 120 148 1408 1172
rect 1472 148 1492 1172
rect 120 120 1492 148
rect -1492 -148 -120 -120
rect -1492 -1172 -204 -148
rect -140 -1172 -120 -148
rect -1492 -1200 -120 -1172
rect 120 -148 1492 -120
rect 120 -1172 1408 -148
rect 1472 -1172 1492 -148
rect 120 -1200 1492 -1172
rect -1492 -1468 -120 -1440
rect -1492 -2492 -204 -1468
rect -140 -2492 -120 -1468
rect -1492 -2520 -120 -2492
rect 120 -1468 1492 -1440
rect 120 -2492 1408 -1468
rect 1472 -2492 1492 -1468
rect 120 -2520 1492 -2492
rect -1492 -2788 -120 -2760
rect -1492 -3812 -204 -2788
rect -140 -3812 -120 -2788
rect -1492 -3840 -120 -3812
rect 120 -2788 1492 -2760
rect 120 -3812 1408 -2788
rect 1472 -3812 1492 -2788
rect 120 -3840 1492 -3812
rect -1492 -4108 -120 -4080
rect -1492 -5132 -204 -4108
rect -140 -5132 -120 -4108
rect -1492 -5160 -120 -5132
rect 120 -4108 1492 -4080
rect 120 -5132 1408 -4108
rect 1472 -5132 1492 -4108
rect 120 -5160 1492 -5132
rect -1492 -5428 -120 -5400
rect -1492 -6452 -204 -5428
rect -140 -6452 -120 -5428
rect -1492 -6480 -120 -6452
rect 120 -5428 1492 -5400
rect 120 -6452 1408 -5428
rect 1472 -6452 1492 -5428
rect 120 -6480 1492 -6452
rect -1492 -6748 -120 -6720
rect -1492 -7772 -204 -6748
rect -140 -7772 -120 -6748
rect -1492 -7800 -120 -7772
rect 120 -6748 1492 -6720
rect 120 -7772 1408 -6748
rect 1472 -7772 1492 -6748
rect 120 -7800 1492 -7772
rect -1492 -8068 -120 -8040
rect -1492 -9092 -204 -8068
rect -140 -9092 -120 -8068
rect -1492 -9120 -120 -9092
rect 120 -8068 1492 -8040
rect 120 -9092 1408 -8068
rect 1472 -9092 1492 -8068
rect 120 -9120 1492 -9092
rect -1492 -9388 -120 -9360
rect -1492 -10412 -204 -9388
rect -140 -10412 -120 -9388
rect -1492 -10440 -120 -10412
rect 120 -9388 1492 -9360
rect 120 -10412 1408 -9388
rect 1472 -10412 1492 -9388
rect 120 -10440 1492 -10412
<< via3 >>
rect -204 9388 -140 10412
rect 1408 9388 1472 10412
rect -204 8068 -140 9092
rect 1408 8068 1472 9092
rect -204 6748 -140 7772
rect 1408 6748 1472 7772
rect -204 5428 -140 6452
rect 1408 5428 1472 6452
rect -204 4108 -140 5132
rect 1408 4108 1472 5132
rect -204 2788 -140 3812
rect 1408 2788 1472 3812
rect -204 1468 -140 2492
rect 1408 1468 1472 2492
rect -204 148 -140 1172
rect 1408 148 1472 1172
rect -204 -1172 -140 -148
rect 1408 -1172 1472 -148
rect -204 -2492 -140 -1468
rect 1408 -2492 1472 -1468
rect -204 -3812 -140 -2788
rect 1408 -3812 1472 -2788
rect -204 -5132 -140 -4108
rect 1408 -5132 1472 -4108
rect -204 -6452 -140 -5428
rect 1408 -6452 1472 -5428
rect -204 -7772 -140 -6748
rect 1408 -7772 1472 -6748
rect -204 -9092 -140 -8068
rect 1408 -9092 1472 -8068
rect -204 -10412 -140 -9388
rect 1408 -10412 1472 -9388
<< mimcap >>
rect -1452 10360 -452 10400
rect -1452 9440 -1412 10360
rect -492 9440 -452 10360
rect -1452 9400 -452 9440
rect 160 10360 1160 10400
rect 160 9440 200 10360
rect 1120 9440 1160 10360
rect 160 9400 1160 9440
rect -1452 9040 -452 9080
rect -1452 8120 -1412 9040
rect -492 8120 -452 9040
rect -1452 8080 -452 8120
rect 160 9040 1160 9080
rect 160 8120 200 9040
rect 1120 8120 1160 9040
rect 160 8080 1160 8120
rect -1452 7720 -452 7760
rect -1452 6800 -1412 7720
rect -492 6800 -452 7720
rect -1452 6760 -452 6800
rect 160 7720 1160 7760
rect 160 6800 200 7720
rect 1120 6800 1160 7720
rect 160 6760 1160 6800
rect -1452 6400 -452 6440
rect -1452 5480 -1412 6400
rect -492 5480 -452 6400
rect -1452 5440 -452 5480
rect 160 6400 1160 6440
rect 160 5480 200 6400
rect 1120 5480 1160 6400
rect 160 5440 1160 5480
rect -1452 5080 -452 5120
rect -1452 4160 -1412 5080
rect -492 4160 -452 5080
rect -1452 4120 -452 4160
rect 160 5080 1160 5120
rect 160 4160 200 5080
rect 1120 4160 1160 5080
rect 160 4120 1160 4160
rect -1452 3760 -452 3800
rect -1452 2840 -1412 3760
rect -492 2840 -452 3760
rect -1452 2800 -452 2840
rect 160 3760 1160 3800
rect 160 2840 200 3760
rect 1120 2840 1160 3760
rect 160 2800 1160 2840
rect -1452 2440 -452 2480
rect -1452 1520 -1412 2440
rect -492 1520 -452 2440
rect -1452 1480 -452 1520
rect 160 2440 1160 2480
rect 160 1520 200 2440
rect 1120 1520 1160 2440
rect 160 1480 1160 1520
rect -1452 1120 -452 1160
rect -1452 200 -1412 1120
rect -492 200 -452 1120
rect -1452 160 -452 200
rect 160 1120 1160 1160
rect 160 200 200 1120
rect 1120 200 1160 1120
rect 160 160 1160 200
rect -1452 -200 -452 -160
rect -1452 -1120 -1412 -200
rect -492 -1120 -452 -200
rect -1452 -1160 -452 -1120
rect 160 -200 1160 -160
rect 160 -1120 200 -200
rect 1120 -1120 1160 -200
rect 160 -1160 1160 -1120
rect -1452 -1520 -452 -1480
rect -1452 -2440 -1412 -1520
rect -492 -2440 -452 -1520
rect -1452 -2480 -452 -2440
rect 160 -1520 1160 -1480
rect 160 -2440 200 -1520
rect 1120 -2440 1160 -1520
rect 160 -2480 1160 -2440
rect -1452 -2840 -452 -2800
rect -1452 -3760 -1412 -2840
rect -492 -3760 -452 -2840
rect -1452 -3800 -452 -3760
rect 160 -2840 1160 -2800
rect 160 -3760 200 -2840
rect 1120 -3760 1160 -2840
rect 160 -3800 1160 -3760
rect -1452 -4160 -452 -4120
rect -1452 -5080 -1412 -4160
rect -492 -5080 -452 -4160
rect -1452 -5120 -452 -5080
rect 160 -4160 1160 -4120
rect 160 -5080 200 -4160
rect 1120 -5080 1160 -4160
rect 160 -5120 1160 -5080
rect -1452 -5480 -452 -5440
rect -1452 -6400 -1412 -5480
rect -492 -6400 -452 -5480
rect -1452 -6440 -452 -6400
rect 160 -5480 1160 -5440
rect 160 -6400 200 -5480
rect 1120 -6400 1160 -5480
rect 160 -6440 1160 -6400
rect -1452 -6800 -452 -6760
rect -1452 -7720 -1412 -6800
rect -492 -7720 -452 -6800
rect -1452 -7760 -452 -7720
rect 160 -6800 1160 -6760
rect 160 -7720 200 -6800
rect 1120 -7720 1160 -6800
rect 160 -7760 1160 -7720
rect -1452 -8120 -452 -8080
rect -1452 -9040 -1412 -8120
rect -492 -9040 -452 -8120
rect -1452 -9080 -452 -9040
rect 160 -8120 1160 -8080
rect 160 -9040 200 -8120
rect 1120 -9040 1160 -8120
rect 160 -9080 1160 -9040
rect -1452 -9440 -452 -9400
rect -1452 -10360 -1412 -9440
rect -492 -10360 -452 -9440
rect -1452 -10400 -452 -10360
rect 160 -9440 1160 -9400
rect 160 -10360 200 -9440
rect 1120 -10360 1160 -9440
rect 160 -10400 1160 -10360
<< mimcapcontact >>
rect -1412 9440 -492 10360
rect 200 9440 1120 10360
rect -1412 8120 -492 9040
rect 200 8120 1120 9040
rect -1412 6800 -492 7720
rect 200 6800 1120 7720
rect -1412 5480 -492 6400
rect 200 5480 1120 6400
rect -1412 4160 -492 5080
rect 200 4160 1120 5080
rect -1412 2840 -492 3760
rect 200 2840 1120 3760
rect -1412 1520 -492 2440
rect 200 1520 1120 2440
rect -1412 200 -492 1120
rect 200 200 1120 1120
rect -1412 -1120 -492 -200
rect 200 -1120 1120 -200
rect -1412 -2440 -492 -1520
rect 200 -2440 1120 -1520
rect -1412 -3760 -492 -2840
rect 200 -3760 1120 -2840
rect -1412 -5080 -492 -4160
rect 200 -5080 1120 -4160
rect -1412 -6400 -492 -5480
rect 200 -6400 1120 -5480
rect -1412 -7720 -492 -6800
rect 200 -7720 1120 -6800
rect -1412 -9040 -492 -8120
rect 200 -9040 1120 -8120
rect -1412 -10360 -492 -9440
rect 200 -10360 1120 -9440
<< metal4 >>
rect -1004 10361 -900 10560
rect -224 10412 -120 10560
rect -1413 10360 -491 10361
rect -1413 9440 -1412 10360
rect -492 9440 -491 10360
rect -1413 9439 -491 9440
rect -1004 9041 -900 9439
rect -224 9388 -204 10412
rect -140 9388 -120 10412
rect 608 10361 712 10560
rect 1388 10412 1492 10560
rect 199 10360 1121 10361
rect 199 9440 200 10360
rect 1120 9440 1121 10360
rect 199 9439 1121 9440
rect -224 9092 -120 9388
rect -1413 9040 -491 9041
rect -1413 8120 -1412 9040
rect -492 8120 -491 9040
rect -1413 8119 -491 8120
rect -1004 7721 -900 8119
rect -224 8068 -204 9092
rect -140 8068 -120 9092
rect 608 9041 712 9439
rect 1388 9388 1408 10412
rect 1472 9388 1492 10412
rect 1388 9092 1492 9388
rect 199 9040 1121 9041
rect 199 8120 200 9040
rect 1120 8120 1121 9040
rect 199 8119 1121 8120
rect -224 7772 -120 8068
rect -1413 7720 -491 7721
rect -1413 6800 -1412 7720
rect -492 6800 -491 7720
rect -1413 6799 -491 6800
rect -1004 6401 -900 6799
rect -224 6748 -204 7772
rect -140 6748 -120 7772
rect 608 7721 712 8119
rect 1388 8068 1408 9092
rect 1472 8068 1492 9092
rect 1388 7772 1492 8068
rect 199 7720 1121 7721
rect 199 6800 200 7720
rect 1120 6800 1121 7720
rect 199 6799 1121 6800
rect -224 6452 -120 6748
rect -1413 6400 -491 6401
rect -1413 5480 -1412 6400
rect -492 5480 -491 6400
rect -1413 5479 -491 5480
rect -1004 5081 -900 5479
rect -224 5428 -204 6452
rect -140 5428 -120 6452
rect 608 6401 712 6799
rect 1388 6748 1408 7772
rect 1472 6748 1492 7772
rect 1388 6452 1492 6748
rect 199 6400 1121 6401
rect 199 5480 200 6400
rect 1120 5480 1121 6400
rect 199 5479 1121 5480
rect -224 5132 -120 5428
rect -1413 5080 -491 5081
rect -1413 4160 -1412 5080
rect -492 4160 -491 5080
rect -1413 4159 -491 4160
rect -1004 3761 -900 4159
rect -224 4108 -204 5132
rect -140 4108 -120 5132
rect 608 5081 712 5479
rect 1388 5428 1408 6452
rect 1472 5428 1492 6452
rect 1388 5132 1492 5428
rect 199 5080 1121 5081
rect 199 4160 200 5080
rect 1120 4160 1121 5080
rect 199 4159 1121 4160
rect -224 3812 -120 4108
rect -1413 3760 -491 3761
rect -1413 2840 -1412 3760
rect -492 2840 -491 3760
rect -1413 2839 -491 2840
rect -1004 2441 -900 2839
rect -224 2788 -204 3812
rect -140 2788 -120 3812
rect 608 3761 712 4159
rect 1388 4108 1408 5132
rect 1472 4108 1492 5132
rect 1388 3812 1492 4108
rect 199 3760 1121 3761
rect 199 2840 200 3760
rect 1120 2840 1121 3760
rect 199 2839 1121 2840
rect -224 2492 -120 2788
rect -1413 2440 -491 2441
rect -1413 1520 -1412 2440
rect -492 1520 -491 2440
rect -1413 1519 -491 1520
rect -1004 1121 -900 1519
rect -224 1468 -204 2492
rect -140 1468 -120 2492
rect 608 2441 712 2839
rect 1388 2788 1408 3812
rect 1472 2788 1492 3812
rect 1388 2492 1492 2788
rect 199 2440 1121 2441
rect 199 1520 200 2440
rect 1120 1520 1121 2440
rect 199 1519 1121 1520
rect -224 1172 -120 1468
rect -1413 1120 -491 1121
rect -1413 200 -1412 1120
rect -492 200 -491 1120
rect -1413 199 -491 200
rect -1004 -199 -900 199
rect -224 148 -204 1172
rect -140 148 -120 1172
rect 608 1121 712 1519
rect 1388 1468 1408 2492
rect 1472 1468 1492 2492
rect 1388 1172 1492 1468
rect 199 1120 1121 1121
rect 199 200 200 1120
rect 1120 200 1121 1120
rect 199 199 1121 200
rect -224 -148 -120 148
rect -1413 -200 -491 -199
rect -1413 -1120 -1412 -200
rect -492 -1120 -491 -200
rect -1413 -1121 -491 -1120
rect -1004 -1519 -900 -1121
rect -224 -1172 -204 -148
rect -140 -1172 -120 -148
rect 608 -199 712 199
rect 1388 148 1408 1172
rect 1472 148 1492 1172
rect 1388 -148 1492 148
rect 199 -200 1121 -199
rect 199 -1120 200 -200
rect 1120 -1120 1121 -200
rect 199 -1121 1121 -1120
rect -224 -1468 -120 -1172
rect -1413 -1520 -491 -1519
rect -1413 -2440 -1412 -1520
rect -492 -2440 -491 -1520
rect -1413 -2441 -491 -2440
rect -1004 -2839 -900 -2441
rect -224 -2492 -204 -1468
rect -140 -2492 -120 -1468
rect 608 -1519 712 -1121
rect 1388 -1172 1408 -148
rect 1472 -1172 1492 -148
rect 1388 -1468 1492 -1172
rect 199 -1520 1121 -1519
rect 199 -2440 200 -1520
rect 1120 -2440 1121 -1520
rect 199 -2441 1121 -2440
rect -224 -2788 -120 -2492
rect -1413 -2840 -491 -2839
rect -1413 -3760 -1412 -2840
rect -492 -3760 -491 -2840
rect -1413 -3761 -491 -3760
rect -1004 -4159 -900 -3761
rect -224 -3812 -204 -2788
rect -140 -3812 -120 -2788
rect 608 -2839 712 -2441
rect 1388 -2492 1408 -1468
rect 1472 -2492 1492 -1468
rect 1388 -2788 1492 -2492
rect 199 -2840 1121 -2839
rect 199 -3760 200 -2840
rect 1120 -3760 1121 -2840
rect 199 -3761 1121 -3760
rect -224 -4108 -120 -3812
rect -1413 -4160 -491 -4159
rect -1413 -5080 -1412 -4160
rect -492 -5080 -491 -4160
rect -1413 -5081 -491 -5080
rect -1004 -5479 -900 -5081
rect -224 -5132 -204 -4108
rect -140 -5132 -120 -4108
rect 608 -4159 712 -3761
rect 1388 -3812 1408 -2788
rect 1472 -3812 1492 -2788
rect 1388 -4108 1492 -3812
rect 199 -4160 1121 -4159
rect 199 -5080 200 -4160
rect 1120 -5080 1121 -4160
rect 199 -5081 1121 -5080
rect -224 -5428 -120 -5132
rect -1413 -5480 -491 -5479
rect -1413 -6400 -1412 -5480
rect -492 -6400 -491 -5480
rect -1413 -6401 -491 -6400
rect -1004 -6799 -900 -6401
rect -224 -6452 -204 -5428
rect -140 -6452 -120 -5428
rect 608 -5479 712 -5081
rect 1388 -5132 1408 -4108
rect 1472 -5132 1492 -4108
rect 1388 -5428 1492 -5132
rect 199 -5480 1121 -5479
rect 199 -6400 200 -5480
rect 1120 -6400 1121 -5480
rect 199 -6401 1121 -6400
rect -224 -6748 -120 -6452
rect -1413 -6800 -491 -6799
rect -1413 -7720 -1412 -6800
rect -492 -7720 -491 -6800
rect -1413 -7721 -491 -7720
rect -1004 -8119 -900 -7721
rect -224 -7772 -204 -6748
rect -140 -7772 -120 -6748
rect 608 -6799 712 -6401
rect 1388 -6452 1408 -5428
rect 1472 -6452 1492 -5428
rect 1388 -6748 1492 -6452
rect 199 -6800 1121 -6799
rect 199 -7720 200 -6800
rect 1120 -7720 1121 -6800
rect 199 -7721 1121 -7720
rect -224 -8068 -120 -7772
rect -1413 -8120 -491 -8119
rect -1413 -9040 -1412 -8120
rect -492 -9040 -491 -8120
rect -1413 -9041 -491 -9040
rect -1004 -9439 -900 -9041
rect -224 -9092 -204 -8068
rect -140 -9092 -120 -8068
rect 608 -8119 712 -7721
rect 1388 -7772 1408 -6748
rect 1472 -7772 1492 -6748
rect 1388 -8068 1492 -7772
rect 199 -8120 1121 -8119
rect 199 -9040 200 -8120
rect 1120 -9040 1121 -8120
rect 199 -9041 1121 -9040
rect -224 -9388 -120 -9092
rect -1413 -9440 -491 -9439
rect -1413 -10360 -1412 -9440
rect -492 -10360 -491 -9440
rect -1413 -10361 -491 -10360
rect -1004 -10560 -900 -10361
rect -224 -10412 -204 -9388
rect -140 -10412 -120 -9388
rect 608 -9439 712 -9041
rect 1388 -9092 1408 -8068
rect 1472 -9092 1492 -8068
rect 1388 -9388 1492 -9092
rect 199 -9440 1121 -9439
rect 199 -10360 200 -9440
rect 1120 -10360 1121 -9440
rect 199 -10361 1121 -10360
rect -224 -10560 -120 -10412
rect 608 -10560 712 -10361
rect 1388 -10412 1408 -9388
rect 1472 -10412 1492 -9388
rect 1388 -10560 1492 -10412
<< properties >>
string FIXED_BBOX 120 9360 1200 10440
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5.0 l 5.0 val 53.8 carea 2.00 cperi 0.19 nx 2 ny 16 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1754800442
<< error_p >>
rect -67 93 -21 105
rect -67 46 -61 93
rect -67 34 -21 46
rect 21 16 67 28
rect 21 -31 27 16
rect 21 -43 67 -31
rect -29 -98 29 -92
rect -29 -132 -17 -98
rect -29 -138 29 -132
<< nmos >>
rect -15 -60 15 122
<< ndiff >>
rect -73 110 -15 122
rect -73 -48 -61 110
rect -27 -48 -15 110
rect -73 -60 -15 -48
rect 15 110 73 122
rect 15 -48 27 110
rect 61 -48 73 110
rect 15 -60 73 -48
<< ndiffc >>
rect -61 -48 -27 110
rect 27 -48 61 110
<< poly >>
rect -15 122 15 148
rect -15 -82 15 -60
rect -33 -98 33 -82
rect -33 -132 -17 -98
rect 17 -132 33 -98
rect -33 -148 33 -132
<< polycont >>
rect -17 -132 17 -98
<< locali >>
rect -61 110 -27 126
rect -61 -64 -27 -48
rect 27 110 61 126
rect 27 -64 61 -48
rect -33 -132 -17 -98
rect 17 -132 33 -98
<< viali >>
rect -61 46 -27 93
rect 27 -31 61 16
rect -17 -132 17 -98
<< metal1 >>
rect -67 93 -21 105
rect -67 46 -61 93
rect -27 46 -21 93
rect -67 34 -21 46
rect 21 16 67 28
rect 21 -31 27 16
rect 61 -31 67 16
rect 21 -43 67 -31
rect -29 -98 29 -92
rect -29 -132 -17 -98
rect 17 -132 29 -98
rect -29 -138 29 -132
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.91 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc +30 viadrn -30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1755037679
<< metal3 >>
rect -6328 5132 -4956 5160
rect -6328 4108 -5040 5132
rect -4976 4108 -4956 5132
rect -6328 4080 -4956 4108
rect -4716 5132 -3344 5160
rect -4716 4108 -3428 5132
rect -3364 4108 -3344 5132
rect -4716 4080 -3344 4108
rect -3104 5132 -1732 5160
rect -3104 4108 -1816 5132
rect -1752 4108 -1732 5132
rect -3104 4080 -1732 4108
rect -1492 5132 -120 5160
rect -1492 4108 -204 5132
rect -140 4108 -120 5132
rect -1492 4080 -120 4108
rect 120 5132 1492 5160
rect 120 4108 1408 5132
rect 1472 4108 1492 5132
rect 120 4080 1492 4108
rect 1732 5132 3104 5160
rect 1732 4108 3020 5132
rect 3084 4108 3104 5132
rect 1732 4080 3104 4108
rect 3344 5132 4716 5160
rect 3344 4108 4632 5132
rect 4696 4108 4716 5132
rect 3344 4080 4716 4108
rect 4956 5132 6328 5160
rect 4956 4108 6244 5132
rect 6308 4108 6328 5132
rect 4956 4080 6328 4108
rect -6328 3812 -4956 3840
rect -6328 2788 -5040 3812
rect -4976 2788 -4956 3812
rect -6328 2760 -4956 2788
rect -4716 3812 -3344 3840
rect -4716 2788 -3428 3812
rect -3364 2788 -3344 3812
rect -4716 2760 -3344 2788
rect -3104 3812 -1732 3840
rect -3104 2788 -1816 3812
rect -1752 2788 -1732 3812
rect -3104 2760 -1732 2788
rect -1492 3812 -120 3840
rect -1492 2788 -204 3812
rect -140 2788 -120 3812
rect -1492 2760 -120 2788
rect 120 3812 1492 3840
rect 120 2788 1408 3812
rect 1472 2788 1492 3812
rect 120 2760 1492 2788
rect 1732 3812 3104 3840
rect 1732 2788 3020 3812
rect 3084 2788 3104 3812
rect 1732 2760 3104 2788
rect 3344 3812 4716 3840
rect 3344 2788 4632 3812
rect 4696 2788 4716 3812
rect 3344 2760 4716 2788
rect 4956 3812 6328 3840
rect 4956 2788 6244 3812
rect 6308 2788 6328 3812
rect 4956 2760 6328 2788
rect -6328 2492 -4956 2520
rect -6328 1468 -5040 2492
rect -4976 1468 -4956 2492
rect -6328 1440 -4956 1468
rect -4716 2492 -3344 2520
rect -4716 1468 -3428 2492
rect -3364 1468 -3344 2492
rect -4716 1440 -3344 1468
rect -3104 2492 -1732 2520
rect -3104 1468 -1816 2492
rect -1752 1468 -1732 2492
rect -3104 1440 -1732 1468
rect -1492 2492 -120 2520
rect -1492 1468 -204 2492
rect -140 1468 -120 2492
rect -1492 1440 -120 1468
rect 120 2492 1492 2520
rect 120 1468 1408 2492
rect 1472 1468 1492 2492
rect 120 1440 1492 1468
rect 1732 2492 3104 2520
rect 1732 1468 3020 2492
rect 3084 1468 3104 2492
rect 1732 1440 3104 1468
rect 3344 2492 4716 2520
rect 3344 1468 4632 2492
rect 4696 1468 4716 2492
rect 3344 1440 4716 1468
rect 4956 2492 6328 2520
rect 4956 1468 6244 2492
rect 6308 1468 6328 2492
rect 4956 1440 6328 1468
rect -6328 1172 -4956 1200
rect -6328 148 -5040 1172
rect -4976 148 -4956 1172
rect -6328 120 -4956 148
rect -4716 1172 -3344 1200
rect -4716 148 -3428 1172
rect -3364 148 -3344 1172
rect -4716 120 -3344 148
rect -3104 1172 -1732 1200
rect -3104 148 -1816 1172
rect -1752 148 -1732 1172
rect -3104 120 -1732 148
rect -1492 1172 -120 1200
rect -1492 148 -204 1172
rect -140 148 -120 1172
rect -1492 120 -120 148
rect 120 1172 1492 1200
rect 120 148 1408 1172
rect 1472 148 1492 1172
rect 120 120 1492 148
rect 1732 1172 3104 1200
rect 1732 148 3020 1172
rect 3084 148 3104 1172
rect 1732 120 3104 148
rect 3344 1172 4716 1200
rect 3344 148 4632 1172
rect 4696 148 4716 1172
rect 3344 120 4716 148
rect 4956 1172 6328 1200
rect 4956 148 6244 1172
rect 6308 148 6328 1172
rect 4956 120 6328 148
rect -6328 -148 -4956 -120
rect -6328 -1172 -5040 -148
rect -4976 -1172 -4956 -148
rect -6328 -1200 -4956 -1172
rect -4716 -148 -3344 -120
rect -4716 -1172 -3428 -148
rect -3364 -1172 -3344 -148
rect -4716 -1200 -3344 -1172
rect -3104 -148 -1732 -120
rect -3104 -1172 -1816 -148
rect -1752 -1172 -1732 -148
rect -3104 -1200 -1732 -1172
rect -1492 -148 -120 -120
rect -1492 -1172 -204 -148
rect -140 -1172 -120 -148
rect -1492 -1200 -120 -1172
rect 120 -148 1492 -120
rect 120 -1172 1408 -148
rect 1472 -1172 1492 -148
rect 120 -1200 1492 -1172
rect 1732 -148 3104 -120
rect 1732 -1172 3020 -148
rect 3084 -1172 3104 -148
rect 1732 -1200 3104 -1172
rect 3344 -148 4716 -120
rect 3344 -1172 4632 -148
rect 4696 -1172 4716 -148
rect 3344 -1200 4716 -1172
rect 4956 -148 6328 -120
rect 4956 -1172 6244 -148
rect 6308 -1172 6328 -148
rect 4956 -1200 6328 -1172
rect -6328 -1468 -4956 -1440
rect -6328 -2492 -5040 -1468
rect -4976 -2492 -4956 -1468
rect -6328 -2520 -4956 -2492
rect -4716 -1468 -3344 -1440
rect -4716 -2492 -3428 -1468
rect -3364 -2492 -3344 -1468
rect -4716 -2520 -3344 -2492
rect -3104 -1468 -1732 -1440
rect -3104 -2492 -1816 -1468
rect -1752 -2492 -1732 -1468
rect -3104 -2520 -1732 -2492
rect -1492 -1468 -120 -1440
rect -1492 -2492 -204 -1468
rect -140 -2492 -120 -1468
rect -1492 -2520 -120 -2492
rect 120 -1468 1492 -1440
rect 120 -2492 1408 -1468
rect 1472 -2492 1492 -1468
rect 120 -2520 1492 -2492
rect 1732 -1468 3104 -1440
rect 1732 -2492 3020 -1468
rect 3084 -2492 3104 -1468
rect 1732 -2520 3104 -2492
rect 3344 -1468 4716 -1440
rect 3344 -2492 4632 -1468
rect 4696 -2492 4716 -1468
rect 3344 -2520 4716 -2492
rect 4956 -1468 6328 -1440
rect 4956 -2492 6244 -1468
rect 6308 -2492 6328 -1468
rect 4956 -2520 6328 -2492
rect -6328 -2788 -4956 -2760
rect -6328 -3812 -5040 -2788
rect -4976 -3812 -4956 -2788
rect -6328 -3840 -4956 -3812
rect -4716 -2788 -3344 -2760
rect -4716 -3812 -3428 -2788
rect -3364 -3812 -3344 -2788
rect -4716 -3840 -3344 -3812
rect -3104 -2788 -1732 -2760
rect -3104 -3812 -1816 -2788
rect -1752 -3812 -1732 -2788
rect -3104 -3840 -1732 -3812
rect -1492 -2788 -120 -2760
rect -1492 -3812 -204 -2788
rect -140 -3812 -120 -2788
rect -1492 -3840 -120 -3812
rect 120 -2788 1492 -2760
rect 120 -3812 1408 -2788
rect 1472 -3812 1492 -2788
rect 120 -3840 1492 -3812
rect 1732 -2788 3104 -2760
rect 1732 -3812 3020 -2788
rect 3084 -3812 3104 -2788
rect 1732 -3840 3104 -3812
rect 3344 -2788 4716 -2760
rect 3344 -3812 4632 -2788
rect 4696 -3812 4716 -2788
rect 3344 -3840 4716 -3812
rect 4956 -2788 6328 -2760
rect 4956 -3812 6244 -2788
rect 6308 -3812 6328 -2788
rect 4956 -3840 6328 -3812
rect -6328 -4108 -4956 -4080
rect -6328 -5132 -5040 -4108
rect -4976 -5132 -4956 -4108
rect -6328 -5160 -4956 -5132
rect -4716 -4108 -3344 -4080
rect -4716 -5132 -3428 -4108
rect -3364 -5132 -3344 -4108
rect -4716 -5160 -3344 -5132
rect -3104 -4108 -1732 -4080
rect -3104 -5132 -1816 -4108
rect -1752 -5132 -1732 -4108
rect -3104 -5160 -1732 -5132
rect -1492 -4108 -120 -4080
rect -1492 -5132 -204 -4108
rect -140 -5132 -120 -4108
rect -1492 -5160 -120 -5132
rect 120 -4108 1492 -4080
rect 120 -5132 1408 -4108
rect 1472 -5132 1492 -4108
rect 120 -5160 1492 -5132
rect 1732 -4108 3104 -4080
rect 1732 -5132 3020 -4108
rect 3084 -5132 3104 -4108
rect 1732 -5160 3104 -5132
rect 3344 -4108 4716 -4080
rect 3344 -5132 4632 -4108
rect 4696 -5132 4716 -4108
rect 3344 -5160 4716 -5132
rect 4956 -4108 6328 -4080
rect 4956 -5132 6244 -4108
rect 6308 -5132 6328 -4108
rect 4956 -5160 6328 -5132
<< via3 >>
rect -5040 4108 -4976 5132
rect -3428 4108 -3364 5132
rect -1816 4108 -1752 5132
rect -204 4108 -140 5132
rect 1408 4108 1472 5132
rect 3020 4108 3084 5132
rect 4632 4108 4696 5132
rect 6244 4108 6308 5132
rect -5040 2788 -4976 3812
rect -3428 2788 -3364 3812
rect -1816 2788 -1752 3812
rect -204 2788 -140 3812
rect 1408 2788 1472 3812
rect 3020 2788 3084 3812
rect 4632 2788 4696 3812
rect 6244 2788 6308 3812
rect -5040 1468 -4976 2492
rect -3428 1468 -3364 2492
rect -1816 1468 -1752 2492
rect -204 1468 -140 2492
rect 1408 1468 1472 2492
rect 3020 1468 3084 2492
rect 4632 1468 4696 2492
rect 6244 1468 6308 2492
rect -5040 148 -4976 1172
rect -3428 148 -3364 1172
rect -1816 148 -1752 1172
rect -204 148 -140 1172
rect 1408 148 1472 1172
rect 3020 148 3084 1172
rect 4632 148 4696 1172
rect 6244 148 6308 1172
rect -5040 -1172 -4976 -148
rect -3428 -1172 -3364 -148
rect -1816 -1172 -1752 -148
rect -204 -1172 -140 -148
rect 1408 -1172 1472 -148
rect 3020 -1172 3084 -148
rect 4632 -1172 4696 -148
rect 6244 -1172 6308 -148
rect -5040 -2492 -4976 -1468
rect -3428 -2492 -3364 -1468
rect -1816 -2492 -1752 -1468
rect -204 -2492 -140 -1468
rect 1408 -2492 1472 -1468
rect 3020 -2492 3084 -1468
rect 4632 -2492 4696 -1468
rect 6244 -2492 6308 -1468
rect -5040 -3812 -4976 -2788
rect -3428 -3812 -3364 -2788
rect -1816 -3812 -1752 -2788
rect -204 -3812 -140 -2788
rect 1408 -3812 1472 -2788
rect 3020 -3812 3084 -2788
rect 4632 -3812 4696 -2788
rect 6244 -3812 6308 -2788
rect -5040 -5132 -4976 -4108
rect -3428 -5132 -3364 -4108
rect -1816 -5132 -1752 -4108
rect -204 -5132 -140 -4108
rect 1408 -5132 1472 -4108
rect 3020 -5132 3084 -4108
rect 4632 -5132 4696 -4108
rect 6244 -5132 6308 -4108
<< mimcap >>
rect -6288 5080 -5288 5120
rect -6288 4160 -6248 5080
rect -5328 4160 -5288 5080
rect -6288 4120 -5288 4160
rect -4676 5080 -3676 5120
rect -4676 4160 -4636 5080
rect -3716 4160 -3676 5080
rect -4676 4120 -3676 4160
rect -3064 5080 -2064 5120
rect -3064 4160 -3024 5080
rect -2104 4160 -2064 5080
rect -3064 4120 -2064 4160
rect -1452 5080 -452 5120
rect -1452 4160 -1412 5080
rect -492 4160 -452 5080
rect -1452 4120 -452 4160
rect 160 5080 1160 5120
rect 160 4160 200 5080
rect 1120 4160 1160 5080
rect 160 4120 1160 4160
rect 1772 5080 2772 5120
rect 1772 4160 1812 5080
rect 2732 4160 2772 5080
rect 1772 4120 2772 4160
rect 3384 5080 4384 5120
rect 3384 4160 3424 5080
rect 4344 4160 4384 5080
rect 3384 4120 4384 4160
rect 4996 5080 5996 5120
rect 4996 4160 5036 5080
rect 5956 4160 5996 5080
rect 4996 4120 5996 4160
rect -6288 3760 -5288 3800
rect -6288 2840 -6248 3760
rect -5328 2840 -5288 3760
rect -6288 2800 -5288 2840
rect -4676 3760 -3676 3800
rect -4676 2840 -4636 3760
rect -3716 2840 -3676 3760
rect -4676 2800 -3676 2840
rect -3064 3760 -2064 3800
rect -3064 2840 -3024 3760
rect -2104 2840 -2064 3760
rect -3064 2800 -2064 2840
rect -1452 3760 -452 3800
rect -1452 2840 -1412 3760
rect -492 2840 -452 3760
rect -1452 2800 -452 2840
rect 160 3760 1160 3800
rect 160 2840 200 3760
rect 1120 2840 1160 3760
rect 160 2800 1160 2840
rect 1772 3760 2772 3800
rect 1772 2840 1812 3760
rect 2732 2840 2772 3760
rect 1772 2800 2772 2840
rect 3384 3760 4384 3800
rect 3384 2840 3424 3760
rect 4344 2840 4384 3760
rect 3384 2800 4384 2840
rect 4996 3760 5996 3800
rect 4996 2840 5036 3760
rect 5956 2840 5996 3760
rect 4996 2800 5996 2840
rect -6288 2440 -5288 2480
rect -6288 1520 -6248 2440
rect -5328 1520 -5288 2440
rect -6288 1480 -5288 1520
rect -4676 2440 -3676 2480
rect -4676 1520 -4636 2440
rect -3716 1520 -3676 2440
rect -4676 1480 -3676 1520
rect -3064 2440 -2064 2480
rect -3064 1520 -3024 2440
rect -2104 1520 -2064 2440
rect -3064 1480 -2064 1520
rect -1452 2440 -452 2480
rect -1452 1520 -1412 2440
rect -492 1520 -452 2440
rect -1452 1480 -452 1520
rect 160 2440 1160 2480
rect 160 1520 200 2440
rect 1120 1520 1160 2440
rect 160 1480 1160 1520
rect 1772 2440 2772 2480
rect 1772 1520 1812 2440
rect 2732 1520 2772 2440
rect 1772 1480 2772 1520
rect 3384 2440 4384 2480
rect 3384 1520 3424 2440
rect 4344 1520 4384 2440
rect 3384 1480 4384 1520
rect 4996 2440 5996 2480
rect 4996 1520 5036 2440
rect 5956 1520 5996 2440
rect 4996 1480 5996 1520
rect -6288 1120 -5288 1160
rect -6288 200 -6248 1120
rect -5328 200 -5288 1120
rect -6288 160 -5288 200
rect -4676 1120 -3676 1160
rect -4676 200 -4636 1120
rect -3716 200 -3676 1120
rect -4676 160 -3676 200
rect -3064 1120 -2064 1160
rect -3064 200 -3024 1120
rect -2104 200 -2064 1120
rect -3064 160 -2064 200
rect -1452 1120 -452 1160
rect -1452 200 -1412 1120
rect -492 200 -452 1120
rect -1452 160 -452 200
rect 160 1120 1160 1160
rect 160 200 200 1120
rect 1120 200 1160 1120
rect 160 160 1160 200
rect 1772 1120 2772 1160
rect 1772 200 1812 1120
rect 2732 200 2772 1120
rect 1772 160 2772 200
rect 3384 1120 4384 1160
rect 3384 200 3424 1120
rect 4344 200 4384 1120
rect 3384 160 4384 200
rect 4996 1120 5996 1160
rect 4996 200 5036 1120
rect 5956 200 5996 1120
rect 4996 160 5996 200
rect -6288 -200 -5288 -160
rect -6288 -1120 -6248 -200
rect -5328 -1120 -5288 -200
rect -6288 -1160 -5288 -1120
rect -4676 -200 -3676 -160
rect -4676 -1120 -4636 -200
rect -3716 -1120 -3676 -200
rect -4676 -1160 -3676 -1120
rect -3064 -200 -2064 -160
rect -3064 -1120 -3024 -200
rect -2104 -1120 -2064 -200
rect -3064 -1160 -2064 -1120
rect -1452 -200 -452 -160
rect -1452 -1120 -1412 -200
rect -492 -1120 -452 -200
rect -1452 -1160 -452 -1120
rect 160 -200 1160 -160
rect 160 -1120 200 -200
rect 1120 -1120 1160 -200
rect 160 -1160 1160 -1120
rect 1772 -200 2772 -160
rect 1772 -1120 1812 -200
rect 2732 -1120 2772 -200
rect 1772 -1160 2772 -1120
rect 3384 -200 4384 -160
rect 3384 -1120 3424 -200
rect 4344 -1120 4384 -200
rect 3384 -1160 4384 -1120
rect 4996 -200 5996 -160
rect 4996 -1120 5036 -200
rect 5956 -1120 5996 -200
rect 4996 -1160 5996 -1120
rect -6288 -1520 -5288 -1480
rect -6288 -2440 -6248 -1520
rect -5328 -2440 -5288 -1520
rect -6288 -2480 -5288 -2440
rect -4676 -1520 -3676 -1480
rect -4676 -2440 -4636 -1520
rect -3716 -2440 -3676 -1520
rect -4676 -2480 -3676 -2440
rect -3064 -1520 -2064 -1480
rect -3064 -2440 -3024 -1520
rect -2104 -2440 -2064 -1520
rect -3064 -2480 -2064 -2440
rect -1452 -1520 -452 -1480
rect -1452 -2440 -1412 -1520
rect -492 -2440 -452 -1520
rect -1452 -2480 -452 -2440
rect 160 -1520 1160 -1480
rect 160 -2440 200 -1520
rect 1120 -2440 1160 -1520
rect 160 -2480 1160 -2440
rect 1772 -1520 2772 -1480
rect 1772 -2440 1812 -1520
rect 2732 -2440 2772 -1520
rect 1772 -2480 2772 -2440
rect 3384 -1520 4384 -1480
rect 3384 -2440 3424 -1520
rect 4344 -2440 4384 -1520
rect 3384 -2480 4384 -2440
rect 4996 -1520 5996 -1480
rect 4996 -2440 5036 -1520
rect 5956 -2440 5996 -1520
rect 4996 -2480 5996 -2440
rect -6288 -2840 -5288 -2800
rect -6288 -3760 -6248 -2840
rect -5328 -3760 -5288 -2840
rect -6288 -3800 -5288 -3760
rect -4676 -2840 -3676 -2800
rect -4676 -3760 -4636 -2840
rect -3716 -3760 -3676 -2840
rect -4676 -3800 -3676 -3760
rect -3064 -2840 -2064 -2800
rect -3064 -3760 -3024 -2840
rect -2104 -3760 -2064 -2840
rect -3064 -3800 -2064 -3760
rect -1452 -2840 -452 -2800
rect -1452 -3760 -1412 -2840
rect -492 -3760 -452 -2840
rect -1452 -3800 -452 -3760
rect 160 -2840 1160 -2800
rect 160 -3760 200 -2840
rect 1120 -3760 1160 -2840
rect 160 -3800 1160 -3760
rect 1772 -2840 2772 -2800
rect 1772 -3760 1812 -2840
rect 2732 -3760 2772 -2840
rect 1772 -3800 2772 -3760
rect 3384 -2840 4384 -2800
rect 3384 -3760 3424 -2840
rect 4344 -3760 4384 -2840
rect 3384 -3800 4384 -3760
rect 4996 -2840 5996 -2800
rect 4996 -3760 5036 -2840
rect 5956 -3760 5996 -2840
rect 4996 -3800 5996 -3760
rect -6288 -4160 -5288 -4120
rect -6288 -5080 -6248 -4160
rect -5328 -5080 -5288 -4160
rect -6288 -5120 -5288 -5080
rect -4676 -4160 -3676 -4120
rect -4676 -5080 -4636 -4160
rect -3716 -5080 -3676 -4160
rect -4676 -5120 -3676 -5080
rect -3064 -4160 -2064 -4120
rect -3064 -5080 -3024 -4160
rect -2104 -5080 -2064 -4160
rect -3064 -5120 -2064 -5080
rect -1452 -4160 -452 -4120
rect -1452 -5080 -1412 -4160
rect -492 -5080 -452 -4160
rect -1452 -5120 -452 -5080
rect 160 -4160 1160 -4120
rect 160 -5080 200 -4160
rect 1120 -5080 1160 -4160
rect 160 -5120 1160 -5080
rect 1772 -4160 2772 -4120
rect 1772 -5080 1812 -4160
rect 2732 -5080 2772 -4160
rect 1772 -5120 2772 -5080
rect 3384 -4160 4384 -4120
rect 3384 -5080 3424 -4160
rect 4344 -5080 4384 -4160
rect 3384 -5120 4384 -5080
rect 4996 -4160 5996 -4120
rect 4996 -5080 5036 -4160
rect 5956 -5080 5996 -4160
rect 4996 -5120 5996 -5080
<< mimcapcontact >>
rect -6248 4160 -5328 5080
rect -4636 4160 -3716 5080
rect -3024 4160 -2104 5080
rect -1412 4160 -492 5080
rect 200 4160 1120 5080
rect 1812 4160 2732 5080
rect 3424 4160 4344 5080
rect 5036 4160 5956 5080
rect -6248 2840 -5328 3760
rect -4636 2840 -3716 3760
rect -3024 2840 -2104 3760
rect -1412 2840 -492 3760
rect 200 2840 1120 3760
rect 1812 2840 2732 3760
rect 3424 2840 4344 3760
rect 5036 2840 5956 3760
rect -6248 1520 -5328 2440
rect -4636 1520 -3716 2440
rect -3024 1520 -2104 2440
rect -1412 1520 -492 2440
rect 200 1520 1120 2440
rect 1812 1520 2732 2440
rect 3424 1520 4344 2440
rect 5036 1520 5956 2440
rect -6248 200 -5328 1120
rect -4636 200 -3716 1120
rect -3024 200 -2104 1120
rect -1412 200 -492 1120
rect 200 200 1120 1120
rect 1812 200 2732 1120
rect 3424 200 4344 1120
rect 5036 200 5956 1120
rect -6248 -1120 -5328 -200
rect -4636 -1120 -3716 -200
rect -3024 -1120 -2104 -200
rect -1412 -1120 -492 -200
rect 200 -1120 1120 -200
rect 1812 -1120 2732 -200
rect 3424 -1120 4344 -200
rect 5036 -1120 5956 -200
rect -6248 -2440 -5328 -1520
rect -4636 -2440 -3716 -1520
rect -3024 -2440 -2104 -1520
rect -1412 -2440 -492 -1520
rect 200 -2440 1120 -1520
rect 1812 -2440 2732 -1520
rect 3424 -2440 4344 -1520
rect 5036 -2440 5956 -1520
rect -6248 -3760 -5328 -2840
rect -4636 -3760 -3716 -2840
rect -3024 -3760 -2104 -2840
rect -1412 -3760 -492 -2840
rect 200 -3760 1120 -2840
rect 1812 -3760 2732 -2840
rect 3424 -3760 4344 -2840
rect 5036 -3760 5956 -2840
rect -6248 -5080 -5328 -4160
rect -4636 -5080 -3716 -4160
rect -3024 -5080 -2104 -4160
rect -1412 -5080 -492 -4160
rect 200 -5080 1120 -4160
rect 1812 -5080 2732 -4160
rect 3424 -5080 4344 -4160
rect 5036 -5080 5956 -4160
<< metal4 >>
rect -5840 5081 -5736 5280
rect -5060 5132 -4956 5280
rect -6249 5080 -5327 5081
rect -6249 4160 -6248 5080
rect -5328 4160 -5327 5080
rect -6249 4159 -5327 4160
rect -5840 3761 -5736 4159
rect -5060 4108 -5040 5132
rect -4976 4108 -4956 5132
rect -4228 5081 -4124 5280
rect -3448 5132 -3344 5280
rect -4637 5080 -3715 5081
rect -4637 4160 -4636 5080
rect -3716 4160 -3715 5080
rect -4637 4159 -3715 4160
rect -5060 3812 -4956 4108
rect -6249 3760 -5327 3761
rect -6249 2840 -6248 3760
rect -5328 2840 -5327 3760
rect -6249 2839 -5327 2840
rect -5840 2441 -5736 2839
rect -5060 2788 -5040 3812
rect -4976 2788 -4956 3812
rect -4228 3761 -4124 4159
rect -3448 4108 -3428 5132
rect -3364 4108 -3344 5132
rect -2616 5081 -2512 5280
rect -1836 5132 -1732 5280
rect -3025 5080 -2103 5081
rect -3025 4160 -3024 5080
rect -2104 4160 -2103 5080
rect -3025 4159 -2103 4160
rect -3448 3812 -3344 4108
rect -4637 3760 -3715 3761
rect -4637 2840 -4636 3760
rect -3716 2840 -3715 3760
rect -4637 2839 -3715 2840
rect -5060 2492 -4956 2788
rect -6249 2440 -5327 2441
rect -6249 1520 -6248 2440
rect -5328 1520 -5327 2440
rect -6249 1519 -5327 1520
rect -5840 1121 -5736 1519
rect -5060 1468 -5040 2492
rect -4976 1468 -4956 2492
rect -4228 2441 -4124 2839
rect -3448 2788 -3428 3812
rect -3364 2788 -3344 3812
rect -2616 3761 -2512 4159
rect -1836 4108 -1816 5132
rect -1752 4108 -1732 5132
rect -1004 5081 -900 5280
rect -224 5132 -120 5280
rect -1413 5080 -491 5081
rect -1413 4160 -1412 5080
rect -492 4160 -491 5080
rect -1413 4159 -491 4160
rect -1836 3812 -1732 4108
rect -3025 3760 -2103 3761
rect -3025 2840 -3024 3760
rect -2104 2840 -2103 3760
rect -3025 2839 -2103 2840
rect -3448 2492 -3344 2788
rect -4637 2440 -3715 2441
rect -4637 1520 -4636 2440
rect -3716 1520 -3715 2440
rect -4637 1519 -3715 1520
rect -5060 1172 -4956 1468
rect -6249 1120 -5327 1121
rect -6249 200 -6248 1120
rect -5328 200 -5327 1120
rect -6249 199 -5327 200
rect -5840 -199 -5736 199
rect -5060 148 -5040 1172
rect -4976 148 -4956 1172
rect -4228 1121 -4124 1519
rect -3448 1468 -3428 2492
rect -3364 1468 -3344 2492
rect -2616 2441 -2512 2839
rect -1836 2788 -1816 3812
rect -1752 2788 -1732 3812
rect -1004 3761 -900 4159
rect -224 4108 -204 5132
rect -140 4108 -120 5132
rect 608 5081 712 5280
rect 1388 5132 1492 5280
rect 199 5080 1121 5081
rect 199 4160 200 5080
rect 1120 4160 1121 5080
rect 199 4159 1121 4160
rect -224 3812 -120 4108
rect -1413 3760 -491 3761
rect -1413 2840 -1412 3760
rect -492 2840 -491 3760
rect -1413 2839 -491 2840
rect -1836 2492 -1732 2788
rect -3025 2440 -2103 2441
rect -3025 1520 -3024 2440
rect -2104 1520 -2103 2440
rect -3025 1519 -2103 1520
rect -3448 1172 -3344 1468
rect -4637 1120 -3715 1121
rect -4637 200 -4636 1120
rect -3716 200 -3715 1120
rect -4637 199 -3715 200
rect -5060 -148 -4956 148
rect -6249 -200 -5327 -199
rect -6249 -1120 -6248 -200
rect -5328 -1120 -5327 -200
rect -6249 -1121 -5327 -1120
rect -5840 -1519 -5736 -1121
rect -5060 -1172 -5040 -148
rect -4976 -1172 -4956 -148
rect -4228 -199 -4124 199
rect -3448 148 -3428 1172
rect -3364 148 -3344 1172
rect -2616 1121 -2512 1519
rect -1836 1468 -1816 2492
rect -1752 1468 -1732 2492
rect -1004 2441 -900 2839
rect -224 2788 -204 3812
rect -140 2788 -120 3812
rect 608 3761 712 4159
rect 1388 4108 1408 5132
rect 1472 4108 1492 5132
rect 2220 5081 2324 5280
rect 3000 5132 3104 5280
rect 1811 5080 2733 5081
rect 1811 4160 1812 5080
rect 2732 4160 2733 5080
rect 1811 4159 2733 4160
rect 1388 3812 1492 4108
rect 199 3760 1121 3761
rect 199 2840 200 3760
rect 1120 2840 1121 3760
rect 199 2839 1121 2840
rect -224 2492 -120 2788
rect -1413 2440 -491 2441
rect -1413 1520 -1412 2440
rect -492 1520 -491 2440
rect -1413 1519 -491 1520
rect -1836 1172 -1732 1468
rect -3025 1120 -2103 1121
rect -3025 200 -3024 1120
rect -2104 200 -2103 1120
rect -3025 199 -2103 200
rect -3448 -148 -3344 148
rect -4637 -200 -3715 -199
rect -4637 -1120 -4636 -200
rect -3716 -1120 -3715 -200
rect -4637 -1121 -3715 -1120
rect -5060 -1468 -4956 -1172
rect -6249 -1520 -5327 -1519
rect -6249 -2440 -6248 -1520
rect -5328 -2440 -5327 -1520
rect -6249 -2441 -5327 -2440
rect -5840 -2839 -5736 -2441
rect -5060 -2492 -5040 -1468
rect -4976 -2492 -4956 -1468
rect -4228 -1519 -4124 -1121
rect -3448 -1172 -3428 -148
rect -3364 -1172 -3344 -148
rect -2616 -199 -2512 199
rect -1836 148 -1816 1172
rect -1752 148 -1732 1172
rect -1004 1121 -900 1519
rect -224 1468 -204 2492
rect -140 1468 -120 2492
rect 608 2441 712 2839
rect 1388 2788 1408 3812
rect 1472 2788 1492 3812
rect 2220 3761 2324 4159
rect 3000 4108 3020 5132
rect 3084 4108 3104 5132
rect 3832 5081 3936 5280
rect 4612 5132 4716 5280
rect 3423 5080 4345 5081
rect 3423 4160 3424 5080
rect 4344 4160 4345 5080
rect 3423 4159 4345 4160
rect 3000 3812 3104 4108
rect 1811 3760 2733 3761
rect 1811 2840 1812 3760
rect 2732 2840 2733 3760
rect 1811 2839 2733 2840
rect 1388 2492 1492 2788
rect 199 2440 1121 2441
rect 199 1520 200 2440
rect 1120 1520 1121 2440
rect 199 1519 1121 1520
rect -224 1172 -120 1468
rect -1413 1120 -491 1121
rect -1413 200 -1412 1120
rect -492 200 -491 1120
rect -1413 199 -491 200
rect -1836 -148 -1732 148
rect -3025 -200 -2103 -199
rect -3025 -1120 -3024 -200
rect -2104 -1120 -2103 -200
rect -3025 -1121 -2103 -1120
rect -3448 -1468 -3344 -1172
rect -4637 -1520 -3715 -1519
rect -4637 -2440 -4636 -1520
rect -3716 -2440 -3715 -1520
rect -4637 -2441 -3715 -2440
rect -5060 -2788 -4956 -2492
rect -6249 -2840 -5327 -2839
rect -6249 -3760 -6248 -2840
rect -5328 -3760 -5327 -2840
rect -6249 -3761 -5327 -3760
rect -5840 -4159 -5736 -3761
rect -5060 -3812 -5040 -2788
rect -4976 -3812 -4956 -2788
rect -4228 -2839 -4124 -2441
rect -3448 -2492 -3428 -1468
rect -3364 -2492 -3344 -1468
rect -2616 -1519 -2512 -1121
rect -1836 -1172 -1816 -148
rect -1752 -1172 -1732 -148
rect -1004 -199 -900 199
rect -224 148 -204 1172
rect -140 148 -120 1172
rect 608 1121 712 1519
rect 1388 1468 1408 2492
rect 1472 1468 1492 2492
rect 2220 2441 2324 2839
rect 3000 2788 3020 3812
rect 3084 2788 3104 3812
rect 3832 3761 3936 4159
rect 4612 4108 4632 5132
rect 4696 4108 4716 5132
rect 5444 5081 5548 5280
rect 6224 5132 6328 5280
rect 5035 5080 5957 5081
rect 5035 4160 5036 5080
rect 5956 4160 5957 5080
rect 5035 4159 5957 4160
rect 4612 3812 4716 4108
rect 3423 3760 4345 3761
rect 3423 2840 3424 3760
rect 4344 2840 4345 3760
rect 3423 2839 4345 2840
rect 3000 2492 3104 2788
rect 1811 2440 2733 2441
rect 1811 1520 1812 2440
rect 2732 1520 2733 2440
rect 1811 1519 2733 1520
rect 1388 1172 1492 1468
rect 199 1120 1121 1121
rect 199 200 200 1120
rect 1120 200 1121 1120
rect 199 199 1121 200
rect -224 -148 -120 148
rect -1413 -200 -491 -199
rect -1413 -1120 -1412 -200
rect -492 -1120 -491 -200
rect -1413 -1121 -491 -1120
rect -1836 -1468 -1732 -1172
rect -3025 -1520 -2103 -1519
rect -3025 -2440 -3024 -1520
rect -2104 -2440 -2103 -1520
rect -3025 -2441 -2103 -2440
rect -3448 -2788 -3344 -2492
rect -4637 -2840 -3715 -2839
rect -4637 -3760 -4636 -2840
rect -3716 -3760 -3715 -2840
rect -4637 -3761 -3715 -3760
rect -5060 -4108 -4956 -3812
rect -6249 -4160 -5327 -4159
rect -6249 -5080 -6248 -4160
rect -5328 -5080 -5327 -4160
rect -6249 -5081 -5327 -5080
rect -5840 -5280 -5736 -5081
rect -5060 -5132 -5040 -4108
rect -4976 -5132 -4956 -4108
rect -4228 -4159 -4124 -3761
rect -3448 -3812 -3428 -2788
rect -3364 -3812 -3344 -2788
rect -2616 -2839 -2512 -2441
rect -1836 -2492 -1816 -1468
rect -1752 -2492 -1732 -1468
rect -1004 -1519 -900 -1121
rect -224 -1172 -204 -148
rect -140 -1172 -120 -148
rect 608 -199 712 199
rect 1388 148 1408 1172
rect 1472 148 1492 1172
rect 2220 1121 2324 1519
rect 3000 1468 3020 2492
rect 3084 1468 3104 2492
rect 3832 2441 3936 2839
rect 4612 2788 4632 3812
rect 4696 2788 4716 3812
rect 5444 3761 5548 4159
rect 6224 4108 6244 5132
rect 6308 4108 6328 5132
rect 6224 3812 6328 4108
rect 5035 3760 5957 3761
rect 5035 2840 5036 3760
rect 5956 2840 5957 3760
rect 5035 2839 5957 2840
rect 4612 2492 4716 2788
rect 3423 2440 4345 2441
rect 3423 1520 3424 2440
rect 4344 1520 4345 2440
rect 3423 1519 4345 1520
rect 3000 1172 3104 1468
rect 1811 1120 2733 1121
rect 1811 200 1812 1120
rect 2732 200 2733 1120
rect 1811 199 2733 200
rect 1388 -148 1492 148
rect 199 -200 1121 -199
rect 199 -1120 200 -200
rect 1120 -1120 1121 -200
rect 199 -1121 1121 -1120
rect -224 -1468 -120 -1172
rect -1413 -1520 -491 -1519
rect -1413 -2440 -1412 -1520
rect -492 -2440 -491 -1520
rect -1413 -2441 -491 -2440
rect -1836 -2788 -1732 -2492
rect -3025 -2840 -2103 -2839
rect -3025 -3760 -3024 -2840
rect -2104 -3760 -2103 -2840
rect -3025 -3761 -2103 -3760
rect -3448 -4108 -3344 -3812
rect -4637 -4160 -3715 -4159
rect -4637 -5080 -4636 -4160
rect -3716 -5080 -3715 -4160
rect -4637 -5081 -3715 -5080
rect -5060 -5280 -4956 -5132
rect -4228 -5280 -4124 -5081
rect -3448 -5132 -3428 -4108
rect -3364 -5132 -3344 -4108
rect -2616 -4159 -2512 -3761
rect -1836 -3812 -1816 -2788
rect -1752 -3812 -1732 -2788
rect -1004 -2839 -900 -2441
rect -224 -2492 -204 -1468
rect -140 -2492 -120 -1468
rect 608 -1519 712 -1121
rect 1388 -1172 1408 -148
rect 1472 -1172 1492 -148
rect 2220 -199 2324 199
rect 3000 148 3020 1172
rect 3084 148 3104 1172
rect 3832 1121 3936 1519
rect 4612 1468 4632 2492
rect 4696 1468 4716 2492
rect 5444 2441 5548 2839
rect 6224 2788 6244 3812
rect 6308 2788 6328 3812
rect 6224 2492 6328 2788
rect 5035 2440 5957 2441
rect 5035 1520 5036 2440
rect 5956 1520 5957 2440
rect 5035 1519 5957 1520
rect 4612 1172 4716 1468
rect 3423 1120 4345 1121
rect 3423 200 3424 1120
rect 4344 200 4345 1120
rect 3423 199 4345 200
rect 3000 -148 3104 148
rect 1811 -200 2733 -199
rect 1811 -1120 1812 -200
rect 2732 -1120 2733 -200
rect 1811 -1121 2733 -1120
rect 1388 -1468 1492 -1172
rect 199 -1520 1121 -1519
rect 199 -2440 200 -1520
rect 1120 -2440 1121 -1520
rect 199 -2441 1121 -2440
rect -224 -2788 -120 -2492
rect -1413 -2840 -491 -2839
rect -1413 -3760 -1412 -2840
rect -492 -3760 -491 -2840
rect -1413 -3761 -491 -3760
rect -1836 -4108 -1732 -3812
rect -3025 -4160 -2103 -4159
rect -3025 -5080 -3024 -4160
rect -2104 -5080 -2103 -4160
rect -3025 -5081 -2103 -5080
rect -3448 -5280 -3344 -5132
rect -2616 -5280 -2512 -5081
rect -1836 -5132 -1816 -4108
rect -1752 -5132 -1732 -4108
rect -1004 -4159 -900 -3761
rect -224 -3812 -204 -2788
rect -140 -3812 -120 -2788
rect 608 -2839 712 -2441
rect 1388 -2492 1408 -1468
rect 1472 -2492 1492 -1468
rect 2220 -1519 2324 -1121
rect 3000 -1172 3020 -148
rect 3084 -1172 3104 -148
rect 3832 -199 3936 199
rect 4612 148 4632 1172
rect 4696 148 4716 1172
rect 5444 1121 5548 1519
rect 6224 1468 6244 2492
rect 6308 1468 6328 2492
rect 6224 1172 6328 1468
rect 5035 1120 5957 1121
rect 5035 200 5036 1120
rect 5956 200 5957 1120
rect 5035 199 5957 200
rect 4612 -148 4716 148
rect 3423 -200 4345 -199
rect 3423 -1120 3424 -200
rect 4344 -1120 4345 -200
rect 3423 -1121 4345 -1120
rect 3000 -1468 3104 -1172
rect 1811 -1520 2733 -1519
rect 1811 -2440 1812 -1520
rect 2732 -2440 2733 -1520
rect 1811 -2441 2733 -2440
rect 1388 -2788 1492 -2492
rect 199 -2840 1121 -2839
rect 199 -3760 200 -2840
rect 1120 -3760 1121 -2840
rect 199 -3761 1121 -3760
rect -224 -4108 -120 -3812
rect -1413 -4160 -491 -4159
rect -1413 -5080 -1412 -4160
rect -492 -5080 -491 -4160
rect -1413 -5081 -491 -5080
rect -1836 -5280 -1732 -5132
rect -1004 -5280 -900 -5081
rect -224 -5132 -204 -4108
rect -140 -5132 -120 -4108
rect 608 -4159 712 -3761
rect 1388 -3812 1408 -2788
rect 1472 -3812 1492 -2788
rect 2220 -2839 2324 -2441
rect 3000 -2492 3020 -1468
rect 3084 -2492 3104 -1468
rect 3832 -1519 3936 -1121
rect 4612 -1172 4632 -148
rect 4696 -1172 4716 -148
rect 5444 -199 5548 199
rect 6224 148 6244 1172
rect 6308 148 6328 1172
rect 6224 -148 6328 148
rect 5035 -200 5957 -199
rect 5035 -1120 5036 -200
rect 5956 -1120 5957 -200
rect 5035 -1121 5957 -1120
rect 4612 -1468 4716 -1172
rect 3423 -1520 4345 -1519
rect 3423 -2440 3424 -1520
rect 4344 -2440 4345 -1520
rect 3423 -2441 4345 -2440
rect 3000 -2788 3104 -2492
rect 1811 -2840 2733 -2839
rect 1811 -3760 1812 -2840
rect 2732 -3760 2733 -2840
rect 1811 -3761 2733 -3760
rect 1388 -4108 1492 -3812
rect 199 -4160 1121 -4159
rect 199 -5080 200 -4160
rect 1120 -5080 1121 -4160
rect 199 -5081 1121 -5080
rect -224 -5280 -120 -5132
rect 608 -5280 712 -5081
rect 1388 -5132 1408 -4108
rect 1472 -5132 1492 -4108
rect 2220 -4159 2324 -3761
rect 3000 -3812 3020 -2788
rect 3084 -3812 3104 -2788
rect 3832 -2839 3936 -2441
rect 4612 -2492 4632 -1468
rect 4696 -2492 4716 -1468
rect 5444 -1519 5548 -1121
rect 6224 -1172 6244 -148
rect 6308 -1172 6328 -148
rect 6224 -1468 6328 -1172
rect 5035 -1520 5957 -1519
rect 5035 -2440 5036 -1520
rect 5956 -2440 5957 -1520
rect 5035 -2441 5957 -2440
rect 4612 -2788 4716 -2492
rect 3423 -2840 4345 -2839
rect 3423 -3760 3424 -2840
rect 4344 -3760 4345 -2840
rect 3423 -3761 4345 -3760
rect 3000 -4108 3104 -3812
rect 1811 -4160 2733 -4159
rect 1811 -5080 1812 -4160
rect 2732 -5080 2733 -4160
rect 1811 -5081 2733 -5080
rect 1388 -5280 1492 -5132
rect 2220 -5280 2324 -5081
rect 3000 -5132 3020 -4108
rect 3084 -5132 3104 -4108
rect 3832 -4159 3936 -3761
rect 4612 -3812 4632 -2788
rect 4696 -3812 4716 -2788
rect 5444 -2839 5548 -2441
rect 6224 -2492 6244 -1468
rect 6308 -2492 6328 -1468
rect 6224 -2788 6328 -2492
rect 5035 -2840 5957 -2839
rect 5035 -3760 5036 -2840
rect 5956 -3760 5957 -2840
rect 5035 -3761 5957 -3760
rect 4612 -4108 4716 -3812
rect 3423 -4160 4345 -4159
rect 3423 -5080 3424 -4160
rect 4344 -5080 4345 -4160
rect 3423 -5081 4345 -5080
rect 3000 -5280 3104 -5132
rect 3832 -5280 3936 -5081
rect 4612 -5132 4632 -4108
rect 4696 -5132 4716 -4108
rect 5444 -4159 5548 -3761
rect 6224 -3812 6244 -2788
rect 6308 -3812 6328 -2788
rect 6224 -4108 6328 -3812
rect 5035 -4160 5957 -4159
rect 5035 -5080 5036 -4160
rect 5956 -5080 5957 -4160
rect 5035 -5081 5957 -5080
rect 4612 -5280 4716 -5132
rect 5444 -5280 5548 -5081
rect 6224 -5132 6244 -4108
rect 6308 -5132 6328 -4108
rect 6224 -5280 6328 -5132
<< properties >>
string FIXED_BBOX 4956 4080 6036 5160
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5 l 5 val 53.8 carea 2.00 cperi 0.19 nx 8 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1754899758
<< metal3 >>
rect -686 20972 686 21000
rect -686 19948 602 20972
rect 666 19948 686 20972
rect -686 19920 686 19948
rect -686 19652 686 19680
rect -686 18628 602 19652
rect 666 18628 686 19652
rect -686 18600 686 18628
rect -686 18332 686 18360
rect -686 17308 602 18332
rect 666 17308 686 18332
rect -686 17280 686 17308
rect -686 17012 686 17040
rect -686 15988 602 17012
rect 666 15988 686 17012
rect -686 15960 686 15988
rect -686 15692 686 15720
rect -686 14668 602 15692
rect 666 14668 686 15692
rect -686 14640 686 14668
rect -686 14372 686 14400
rect -686 13348 602 14372
rect 666 13348 686 14372
rect -686 13320 686 13348
rect -686 13052 686 13080
rect -686 12028 602 13052
rect 666 12028 686 13052
rect -686 12000 686 12028
rect -686 11732 686 11760
rect -686 10708 602 11732
rect 666 10708 686 11732
rect -686 10680 686 10708
rect -686 10412 686 10440
rect -686 9388 602 10412
rect 666 9388 686 10412
rect -686 9360 686 9388
rect -686 9092 686 9120
rect -686 8068 602 9092
rect 666 8068 686 9092
rect -686 8040 686 8068
rect -686 7772 686 7800
rect -686 6748 602 7772
rect 666 6748 686 7772
rect -686 6720 686 6748
rect -686 6452 686 6480
rect -686 5428 602 6452
rect 666 5428 686 6452
rect -686 5400 686 5428
rect -686 5132 686 5160
rect -686 4108 602 5132
rect 666 4108 686 5132
rect -686 4080 686 4108
rect -686 3812 686 3840
rect -686 2788 602 3812
rect 666 2788 686 3812
rect -686 2760 686 2788
rect -686 2492 686 2520
rect -686 1468 602 2492
rect 666 1468 686 2492
rect -686 1440 686 1468
rect -686 1172 686 1200
rect -686 148 602 1172
rect 666 148 686 1172
rect -686 120 686 148
rect -686 -148 686 -120
rect -686 -1172 602 -148
rect 666 -1172 686 -148
rect -686 -1200 686 -1172
rect -686 -1468 686 -1440
rect -686 -2492 602 -1468
rect 666 -2492 686 -1468
rect -686 -2520 686 -2492
rect -686 -2788 686 -2760
rect -686 -3812 602 -2788
rect 666 -3812 686 -2788
rect -686 -3840 686 -3812
rect -686 -4108 686 -4080
rect -686 -5132 602 -4108
rect 666 -5132 686 -4108
rect -686 -5160 686 -5132
rect -686 -5428 686 -5400
rect -686 -6452 602 -5428
rect 666 -6452 686 -5428
rect -686 -6480 686 -6452
rect -686 -6748 686 -6720
rect -686 -7772 602 -6748
rect 666 -7772 686 -6748
rect -686 -7800 686 -7772
rect -686 -8068 686 -8040
rect -686 -9092 602 -8068
rect 666 -9092 686 -8068
rect -686 -9120 686 -9092
rect -686 -9388 686 -9360
rect -686 -10412 602 -9388
rect 666 -10412 686 -9388
rect -686 -10440 686 -10412
rect -686 -10708 686 -10680
rect -686 -11732 602 -10708
rect 666 -11732 686 -10708
rect -686 -11760 686 -11732
rect -686 -12028 686 -12000
rect -686 -13052 602 -12028
rect 666 -13052 686 -12028
rect -686 -13080 686 -13052
rect -686 -13348 686 -13320
rect -686 -14372 602 -13348
rect 666 -14372 686 -13348
rect -686 -14400 686 -14372
rect -686 -14668 686 -14640
rect -686 -15692 602 -14668
rect 666 -15692 686 -14668
rect -686 -15720 686 -15692
rect -686 -15988 686 -15960
rect -686 -17012 602 -15988
rect 666 -17012 686 -15988
rect -686 -17040 686 -17012
rect -686 -17308 686 -17280
rect -686 -18332 602 -17308
rect 666 -18332 686 -17308
rect -686 -18360 686 -18332
rect -686 -18628 686 -18600
rect -686 -19652 602 -18628
rect 666 -19652 686 -18628
rect -686 -19680 686 -19652
rect -686 -19948 686 -19920
rect -686 -20972 602 -19948
rect 666 -20972 686 -19948
rect -686 -21000 686 -20972
<< via3 >>
rect 602 19948 666 20972
rect 602 18628 666 19652
rect 602 17308 666 18332
rect 602 15988 666 17012
rect 602 14668 666 15692
rect 602 13348 666 14372
rect 602 12028 666 13052
rect 602 10708 666 11732
rect 602 9388 666 10412
rect 602 8068 666 9092
rect 602 6748 666 7772
rect 602 5428 666 6452
rect 602 4108 666 5132
rect 602 2788 666 3812
rect 602 1468 666 2492
rect 602 148 666 1172
rect 602 -1172 666 -148
rect 602 -2492 666 -1468
rect 602 -3812 666 -2788
rect 602 -5132 666 -4108
rect 602 -6452 666 -5428
rect 602 -7772 666 -6748
rect 602 -9092 666 -8068
rect 602 -10412 666 -9388
rect 602 -11732 666 -10708
rect 602 -13052 666 -12028
rect 602 -14372 666 -13348
rect 602 -15692 666 -14668
rect 602 -17012 666 -15988
rect 602 -18332 666 -17308
rect 602 -19652 666 -18628
rect 602 -20972 666 -19948
<< mimcap >>
rect -646 20920 354 20960
rect -646 20000 -606 20920
rect 314 20000 354 20920
rect -646 19960 354 20000
rect -646 19600 354 19640
rect -646 18680 -606 19600
rect 314 18680 354 19600
rect -646 18640 354 18680
rect -646 18280 354 18320
rect -646 17360 -606 18280
rect 314 17360 354 18280
rect -646 17320 354 17360
rect -646 16960 354 17000
rect -646 16040 -606 16960
rect 314 16040 354 16960
rect -646 16000 354 16040
rect -646 15640 354 15680
rect -646 14720 -606 15640
rect 314 14720 354 15640
rect -646 14680 354 14720
rect -646 14320 354 14360
rect -646 13400 -606 14320
rect 314 13400 354 14320
rect -646 13360 354 13400
rect -646 13000 354 13040
rect -646 12080 -606 13000
rect 314 12080 354 13000
rect -646 12040 354 12080
rect -646 11680 354 11720
rect -646 10760 -606 11680
rect 314 10760 354 11680
rect -646 10720 354 10760
rect -646 10360 354 10400
rect -646 9440 -606 10360
rect 314 9440 354 10360
rect -646 9400 354 9440
rect -646 9040 354 9080
rect -646 8120 -606 9040
rect 314 8120 354 9040
rect -646 8080 354 8120
rect -646 7720 354 7760
rect -646 6800 -606 7720
rect 314 6800 354 7720
rect -646 6760 354 6800
rect -646 6400 354 6440
rect -646 5480 -606 6400
rect 314 5480 354 6400
rect -646 5440 354 5480
rect -646 5080 354 5120
rect -646 4160 -606 5080
rect 314 4160 354 5080
rect -646 4120 354 4160
rect -646 3760 354 3800
rect -646 2840 -606 3760
rect 314 2840 354 3760
rect -646 2800 354 2840
rect -646 2440 354 2480
rect -646 1520 -606 2440
rect 314 1520 354 2440
rect -646 1480 354 1520
rect -646 1120 354 1160
rect -646 200 -606 1120
rect 314 200 354 1120
rect -646 160 354 200
rect -646 -200 354 -160
rect -646 -1120 -606 -200
rect 314 -1120 354 -200
rect -646 -1160 354 -1120
rect -646 -1520 354 -1480
rect -646 -2440 -606 -1520
rect 314 -2440 354 -1520
rect -646 -2480 354 -2440
rect -646 -2840 354 -2800
rect -646 -3760 -606 -2840
rect 314 -3760 354 -2840
rect -646 -3800 354 -3760
rect -646 -4160 354 -4120
rect -646 -5080 -606 -4160
rect 314 -5080 354 -4160
rect -646 -5120 354 -5080
rect -646 -5480 354 -5440
rect -646 -6400 -606 -5480
rect 314 -6400 354 -5480
rect -646 -6440 354 -6400
rect -646 -6800 354 -6760
rect -646 -7720 -606 -6800
rect 314 -7720 354 -6800
rect -646 -7760 354 -7720
rect -646 -8120 354 -8080
rect -646 -9040 -606 -8120
rect 314 -9040 354 -8120
rect -646 -9080 354 -9040
rect -646 -9440 354 -9400
rect -646 -10360 -606 -9440
rect 314 -10360 354 -9440
rect -646 -10400 354 -10360
rect -646 -10760 354 -10720
rect -646 -11680 -606 -10760
rect 314 -11680 354 -10760
rect -646 -11720 354 -11680
rect -646 -12080 354 -12040
rect -646 -13000 -606 -12080
rect 314 -13000 354 -12080
rect -646 -13040 354 -13000
rect -646 -13400 354 -13360
rect -646 -14320 -606 -13400
rect 314 -14320 354 -13400
rect -646 -14360 354 -14320
rect -646 -14720 354 -14680
rect -646 -15640 -606 -14720
rect 314 -15640 354 -14720
rect -646 -15680 354 -15640
rect -646 -16040 354 -16000
rect -646 -16960 -606 -16040
rect 314 -16960 354 -16040
rect -646 -17000 354 -16960
rect -646 -17360 354 -17320
rect -646 -18280 -606 -17360
rect 314 -18280 354 -17360
rect -646 -18320 354 -18280
rect -646 -18680 354 -18640
rect -646 -19600 -606 -18680
rect 314 -19600 354 -18680
rect -646 -19640 354 -19600
rect -646 -20000 354 -19960
rect -646 -20920 -606 -20000
rect 314 -20920 354 -20000
rect -646 -20960 354 -20920
<< mimcapcontact >>
rect -606 20000 314 20920
rect -606 18680 314 19600
rect -606 17360 314 18280
rect -606 16040 314 16960
rect -606 14720 314 15640
rect -606 13400 314 14320
rect -606 12080 314 13000
rect -606 10760 314 11680
rect -606 9440 314 10360
rect -606 8120 314 9040
rect -606 6800 314 7720
rect -606 5480 314 6400
rect -606 4160 314 5080
rect -606 2840 314 3760
rect -606 1520 314 2440
rect -606 200 314 1120
rect -606 -1120 314 -200
rect -606 -2440 314 -1520
rect -606 -3760 314 -2840
rect -606 -5080 314 -4160
rect -606 -6400 314 -5480
rect -606 -7720 314 -6800
rect -606 -9040 314 -8120
rect -606 -10360 314 -9440
rect -606 -11680 314 -10760
rect -606 -13000 314 -12080
rect -606 -14320 314 -13400
rect -606 -15640 314 -14720
rect -606 -16960 314 -16040
rect -606 -18280 314 -17360
rect -606 -19600 314 -18680
rect -606 -20920 314 -20000
<< metal4 >>
rect -198 20921 -94 21120
rect 582 20972 686 21120
rect -607 20920 315 20921
rect -607 20000 -606 20920
rect 314 20000 315 20920
rect -607 19999 315 20000
rect -198 19601 -94 19999
rect 582 19948 602 20972
rect 666 19948 686 20972
rect 582 19652 686 19948
rect -607 19600 315 19601
rect -607 18680 -606 19600
rect 314 18680 315 19600
rect -607 18679 315 18680
rect -198 18281 -94 18679
rect 582 18628 602 19652
rect 666 18628 686 19652
rect 582 18332 686 18628
rect -607 18280 315 18281
rect -607 17360 -606 18280
rect 314 17360 315 18280
rect -607 17359 315 17360
rect -198 16961 -94 17359
rect 582 17308 602 18332
rect 666 17308 686 18332
rect 582 17012 686 17308
rect -607 16960 315 16961
rect -607 16040 -606 16960
rect 314 16040 315 16960
rect -607 16039 315 16040
rect -198 15641 -94 16039
rect 582 15988 602 17012
rect 666 15988 686 17012
rect 582 15692 686 15988
rect -607 15640 315 15641
rect -607 14720 -606 15640
rect 314 14720 315 15640
rect -607 14719 315 14720
rect -198 14321 -94 14719
rect 582 14668 602 15692
rect 666 14668 686 15692
rect 582 14372 686 14668
rect -607 14320 315 14321
rect -607 13400 -606 14320
rect 314 13400 315 14320
rect -607 13399 315 13400
rect -198 13001 -94 13399
rect 582 13348 602 14372
rect 666 13348 686 14372
rect 582 13052 686 13348
rect -607 13000 315 13001
rect -607 12080 -606 13000
rect 314 12080 315 13000
rect -607 12079 315 12080
rect -198 11681 -94 12079
rect 582 12028 602 13052
rect 666 12028 686 13052
rect 582 11732 686 12028
rect -607 11680 315 11681
rect -607 10760 -606 11680
rect 314 10760 315 11680
rect -607 10759 315 10760
rect -198 10361 -94 10759
rect 582 10708 602 11732
rect 666 10708 686 11732
rect 582 10412 686 10708
rect -607 10360 315 10361
rect -607 9440 -606 10360
rect 314 9440 315 10360
rect -607 9439 315 9440
rect -198 9041 -94 9439
rect 582 9388 602 10412
rect 666 9388 686 10412
rect 582 9092 686 9388
rect -607 9040 315 9041
rect -607 8120 -606 9040
rect 314 8120 315 9040
rect -607 8119 315 8120
rect -198 7721 -94 8119
rect 582 8068 602 9092
rect 666 8068 686 9092
rect 582 7772 686 8068
rect -607 7720 315 7721
rect -607 6800 -606 7720
rect 314 6800 315 7720
rect -607 6799 315 6800
rect -198 6401 -94 6799
rect 582 6748 602 7772
rect 666 6748 686 7772
rect 582 6452 686 6748
rect -607 6400 315 6401
rect -607 5480 -606 6400
rect 314 5480 315 6400
rect -607 5479 315 5480
rect -198 5081 -94 5479
rect 582 5428 602 6452
rect 666 5428 686 6452
rect 582 5132 686 5428
rect -607 5080 315 5081
rect -607 4160 -606 5080
rect 314 4160 315 5080
rect -607 4159 315 4160
rect -198 3761 -94 4159
rect 582 4108 602 5132
rect 666 4108 686 5132
rect 582 3812 686 4108
rect -607 3760 315 3761
rect -607 2840 -606 3760
rect 314 2840 315 3760
rect -607 2839 315 2840
rect -198 2441 -94 2839
rect 582 2788 602 3812
rect 666 2788 686 3812
rect 582 2492 686 2788
rect -607 2440 315 2441
rect -607 1520 -606 2440
rect 314 1520 315 2440
rect -607 1519 315 1520
rect -198 1121 -94 1519
rect 582 1468 602 2492
rect 666 1468 686 2492
rect 582 1172 686 1468
rect -607 1120 315 1121
rect -607 200 -606 1120
rect 314 200 315 1120
rect -607 199 315 200
rect -198 -199 -94 199
rect 582 148 602 1172
rect 666 148 686 1172
rect 582 -148 686 148
rect -607 -200 315 -199
rect -607 -1120 -606 -200
rect 314 -1120 315 -200
rect -607 -1121 315 -1120
rect -198 -1519 -94 -1121
rect 582 -1172 602 -148
rect 666 -1172 686 -148
rect 582 -1468 686 -1172
rect -607 -1520 315 -1519
rect -607 -2440 -606 -1520
rect 314 -2440 315 -1520
rect -607 -2441 315 -2440
rect -198 -2839 -94 -2441
rect 582 -2492 602 -1468
rect 666 -2492 686 -1468
rect 582 -2788 686 -2492
rect -607 -2840 315 -2839
rect -607 -3760 -606 -2840
rect 314 -3760 315 -2840
rect -607 -3761 315 -3760
rect -198 -4159 -94 -3761
rect 582 -3812 602 -2788
rect 666 -3812 686 -2788
rect 582 -4108 686 -3812
rect -607 -4160 315 -4159
rect -607 -5080 -606 -4160
rect 314 -5080 315 -4160
rect -607 -5081 315 -5080
rect -198 -5479 -94 -5081
rect 582 -5132 602 -4108
rect 666 -5132 686 -4108
rect 582 -5428 686 -5132
rect -607 -5480 315 -5479
rect -607 -6400 -606 -5480
rect 314 -6400 315 -5480
rect -607 -6401 315 -6400
rect -198 -6799 -94 -6401
rect 582 -6452 602 -5428
rect 666 -6452 686 -5428
rect 582 -6748 686 -6452
rect -607 -6800 315 -6799
rect -607 -7720 -606 -6800
rect 314 -7720 315 -6800
rect -607 -7721 315 -7720
rect -198 -8119 -94 -7721
rect 582 -7772 602 -6748
rect 666 -7772 686 -6748
rect 582 -8068 686 -7772
rect -607 -8120 315 -8119
rect -607 -9040 -606 -8120
rect 314 -9040 315 -8120
rect -607 -9041 315 -9040
rect -198 -9439 -94 -9041
rect 582 -9092 602 -8068
rect 666 -9092 686 -8068
rect 582 -9388 686 -9092
rect -607 -9440 315 -9439
rect -607 -10360 -606 -9440
rect 314 -10360 315 -9440
rect -607 -10361 315 -10360
rect -198 -10759 -94 -10361
rect 582 -10412 602 -9388
rect 666 -10412 686 -9388
rect 582 -10708 686 -10412
rect -607 -10760 315 -10759
rect -607 -11680 -606 -10760
rect 314 -11680 315 -10760
rect -607 -11681 315 -11680
rect -198 -12079 -94 -11681
rect 582 -11732 602 -10708
rect 666 -11732 686 -10708
rect 582 -12028 686 -11732
rect -607 -12080 315 -12079
rect -607 -13000 -606 -12080
rect 314 -13000 315 -12080
rect -607 -13001 315 -13000
rect -198 -13399 -94 -13001
rect 582 -13052 602 -12028
rect 666 -13052 686 -12028
rect 582 -13348 686 -13052
rect -607 -13400 315 -13399
rect -607 -14320 -606 -13400
rect 314 -14320 315 -13400
rect -607 -14321 315 -14320
rect -198 -14719 -94 -14321
rect 582 -14372 602 -13348
rect 666 -14372 686 -13348
rect 582 -14668 686 -14372
rect -607 -14720 315 -14719
rect -607 -15640 -606 -14720
rect 314 -15640 315 -14720
rect -607 -15641 315 -15640
rect -198 -16039 -94 -15641
rect 582 -15692 602 -14668
rect 666 -15692 686 -14668
rect 582 -15988 686 -15692
rect -607 -16040 315 -16039
rect -607 -16960 -606 -16040
rect 314 -16960 315 -16040
rect -607 -16961 315 -16960
rect -198 -17359 -94 -16961
rect 582 -17012 602 -15988
rect 666 -17012 686 -15988
rect 582 -17308 686 -17012
rect -607 -17360 315 -17359
rect -607 -18280 -606 -17360
rect 314 -18280 315 -17360
rect -607 -18281 315 -18280
rect -198 -18679 -94 -18281
rect 582 -18332 602 -17308
rect 666 -18332 686 -17308
rect 582 -18628 686 -18332
rect -607 -18680 315 -18679
rect -607 -19600 -606 -18680
rect 314 -19600 315 -18680
rect -607 -19601 315 -19600
rect -198 -19999 -94 -19601
rect 582 -19652 602 -18628
rect 666 -19652 686 -18628
rect 582 -19948 686 -19652
rect -607 -20000 315 -19999
rect -607 -20920 -606 -20000
rect 314 -20920 315 -20000
rect -607 -20921 315 -20920
rect -198 -21120 -94 -20921
rect 582 -20972 602 -19948
rect 666 -20972 686 -19948
rect 582 -21120 686 -20972
<< properties >>
string FIXED_BBOX -686 19920 394 21000
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5.0 l 5.0 val 53.8 carea 2.00 cperi 0.19 nx 1 ny 32 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1754255629
<< error_p >>
rect -29 163 29 169
rect -29 129 -17 163
rect -29 123 29 129
rect -29 -129 29 -123
rect -29 -163 -17 -129
rect -29 -169 29 -163
<< pwell >>
rect -211 -301 211 301
<< nmos >>
rect -15 -91 15 91
<< ndiff >>
rect -73 79 -15 91
rect -73 -79 -61 79
rect -27 -79 -15 79
rect -73 -91 -15 -79
rect 15 79 73 91
rect 15 -79 27 79
rect 61 -79 73 79
rect 15 -91 73 -79
<< ndiffc >>
rect -61 -79 -27 79
rect 27 -79 61 79
<< psubdiff >>
rect -175 231 -79 265
rect 79 231 175 265
rect -175 169 -141 231
rect 141 169 175 231
rect -175 -231 -141 -169
rect 141 -231 175 -169
rect -175 -265 -79 -231
rect 79 -265 175 -231
<< psubdiffcont >>
rect -79 231 79 265
rect -175 -169 -141 169
rect 141 -169 175 169
rect -79 -265 79 -231
<< poly >>
rect -33 163 33 179
rect -33 129 -17 163
rect 17 129 33 163
rect -33 113 33 129
rect -15 91 15 113
rect -15 -113 15 -91
rect -33 -129 33 -113
rect -33 -163 -17 -129
rect 17 -163 33 -129
rect -33 -179 33 -163
<< polycont >>
rect -17 129 17 163
rect -17 -163 17 -129
<< locali >>
rect -175 231 -79 265
rect 79 231 175 265
rect -175 169 -141 231
rect 141 169 175 231
rect -33 129 -17 163
rect 17 129 33 163
rect -61 79 -27 95
rect -61 -95 -27 -79
rect 27 79 61 95
rect 27 -95 61 -79
rect -33 -163 -17 -129
rect 17 -163 33 -129
rect -175 -231 -141 -169
rect 141 -231 175 -169
rect -175 -265 -79 -231
rect 79 -265 175 -231
<< viali >>
rect -17 129 17 163
rect -61 -79 -27 79
rect 27 -79 61 79
rect -17 -163 17 -129
<< metal1 >>
rect -29 163 29 169
rect -29 129 -17 163
rect 17 129 29 163
rect -29 123 29 129
rect -67 79 -21 91
rect -67 -79 -61 79
rect -27 -79 -21 79
rect -67 -91 -21 -79
rect 21 79 67 91
rect 21 -79 27 79
rect 61 -79 67 79
rect 21 -91 67 -79
rect -29 -129 29 -123
rect -29 -163 -17 -129
rect 17 -163 29 -129
rect -29 -169 29 -163
<< properties >>
string FIXED_BBOX -158 -248 158 248
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.91 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

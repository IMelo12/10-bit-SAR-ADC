VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO digital
  CLASS BLOCK ;
  FOREIGN digital ;
  ORIGIN 0.000 0.000 ;
  SIZE 109.400 BY 120.120 ;
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END VDD
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 29.210 10.640 30.810 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.705 10.640 55.305 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.200 10.640 79.800 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 102.695 10.640 104.295 109.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 16.965 10.640 18.565 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.460 10.640 43.060 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 65.955 10.640 67.555 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 90.450 10.640 92.050 109.040 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 105.400 99.320 109.400 99.920 ;
    END
  END clk
  PIN clr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 105.400 107.480 109.400 108.080 ;
    END
  END clr
  PIN comp_clk
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END comp_clk
  PIN comp_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END comp_n
  PIN comp_p
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END comp_p
  PIN done
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 105.400 91.160 109.400 91.760 ;
    END
  END done
  PIN obit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 105.400 83.000 109.400 83.600 ;
    END
  END obit1
  PIN obit10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 105.400 9.560 109.400 10.160 ;
    END
  END obit10
  PIN obit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 105.400 74.840 109.400 75.440 ;
    END
  END obit2
  PIN obit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 105.400 66.680 109.400 67.280 ;
    END
  END obit3
  PIN obit4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 105.400 58.520 109.400 59.120 ;
    END
  END obit4
  PIN obit5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 105.400 50.360 109.400 50.960 ;
    END
  END obit5
  PIN obit6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 105.400 42.200 109.400 42.800 ;
    END
  END obit6
  PIN obit7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 105.400 34.040 109.400 34.640 ;
    END
  END obit7
  PIN obit8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 105.400 25.880 109.400 26.480 ;
    END
  END obit8
  PIN obit9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 105.400 17.720 109.400 18.320 ;
    END
  END obit9
  PIN sw_n1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END sw_n1
  PIN sw_n2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END sw_n2
  PIN sw_n3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END sw_n3
  PIN sw_n4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END sw_n4
  PIN sw_n5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END sw_n5
  PIN sw_n6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END sw_n6
  PIN sw_n7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END sw_n7
  PIN sw_n8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END sw_n8
  PIN sw_n_sp1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END sw_n_sp1
  PIN sw_n_sp2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END sw_n_sp2
  PIN sw_n_sp3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END sw_n_sp3
  PIN sw_n_sp4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END sw_n_sp4
  PIN sw_n_sp5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END sw_n_sp5
  PIN sw_n_sp6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END sw_n_sp6
  PIN sw_n_sp7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END sw_n_sp7
  PIN sw_n_sp8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END sw_n_sp8
  PIN sw_n_sp9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END sw_n_sp9
  PIN sw_p1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 93.010 116.120 93.290 120.120 ;
    END
  END sw_p1
  PIN sw_p2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 86.570 116.120 86.850 120.120 ;
    END
  END sw_p2
  PIN sw_p3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 60.810 116.120 61.090 120.120 ;
    END
  END sw_p3
  PIN sw_p4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.370 116.120 54.650 120.120 ;
    END
  END sw_p4
  PIN sw_p5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 47.930 116.120 48.210 120.120 ;
    END
  END sw_p5
  PIN sw_p6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 22.170 116.120 22.450 120.120 ;
    END
  END sw_p6
  PIN sw_p7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 15.730 116.120 16.010 120.120 ;
    END
  END sw_p7
  PIN sw_p8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 9.290 116.120 9.570 120.120 ;
    END
  END sw_p8
  PIN sw_p_sp1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 105.890 116.120 106.170 120.120 ;
    END
  END sw_p_sp1
  PIN sw_p_sp2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 99.450 116.120 99.730 120.120 ;
    END
  END sw_p_sp2
  PIN sw_p_sp3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 80.130 116.120 80.410 120.120 ;
    END
  END sw_p_sp3
  PIN sw_p_sp4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 73.690 116.120 73.970 120.120 ;
    END
  END sw_p_sp4
  PIN sw_p_sp5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 67.250 116.120 67.530 120.120 ;
    END
  END sw_p_sp5
  PIN sw_p_sp6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 41.490 116.120 41.770 120.120 ;
    END
  END sw_p_sp6
  PIN sw_p_sp7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.050 116.120 35.330 120.120 ;
    END
  END sw_p_sp7
  PIN sw_p_sp8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 28.610 116.120 28.890 120.120 ;
    END
  END sw_p_sp8
  PIN sw_p_sp9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 2.850 116.120 3.130 120.120 ;
    END
  END sw_p_sp9
  PIN sw_sample
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END sw_sample
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 103.500 108.885 ;
      LAYER met1 ;
        RECT 2.830 10.640 106.190 109.040 ;
      LAYER met2 ;
        RECT 3.410 115.840 9.010 116.690 ;
        RECT 9.850 115.840 15.450 116.690 ;
        RECT 16.290 115.840 21.890 116.690 ;
        RECT 22.730 115.840 28.330 116.690 ;
        RECT 29.170 115.840 34.770 116.690 ;
        RECT 35.610 115.840 41.210 116.690 ;
        RECT 42.050 115.840 47.650 116.690 ;
        RECT 48.490 115.840 54.090 116.690 ;
        RECT 54.930 115.840 60.530 116.690 ;
        RECT 61.370 115.840 66.970 116.690 ;
        RECT 67.810 115.840 73.410 116.690 ;
        RECT 74.250 115.840 79.850 116.690 ;
        RECT 80.690 115.840 86.290 116.690 ;
        RECT 87.130 115.840 92.730 116.690 ;
        RECT 93.570 115.840 99.170 116.690 ;
        RECT 100.010 115.840 105.610 116.690 ;
        RECT 2.860 4.280 106.160 115.840 ;
        RECT 3.410 3.670 9.010 4.280 ;
        RECT 9.850 3.670 15.450 4.280 ;
        RECT 16.290 3.670 21.890 4.280 ;
        RECT 22.730 3.670 28.330 4.280 ;
        RECT 29.170 3.670 34.770 4.280 ;
        RECT 35.610 3.670 41.210 4.280 ;
        RECT 42.050 3.670 47.650 4.280 ;
        RECT 48.490 3.670 54.090 4.280 ;
        RECT 54.930 3.670 60.530 4.280 ;
        RECT 61.370 3.670 66.970 4.280 ;
        RECT 67.810 3.670 73.410 4.280 ;
        RECT 74.250 3.670 79.850 4.280 ;
        RECT 80.690 3.670 86.290 4.280 ;
        RECT 87.130 3.670 92.730 4.280 ;
        RECT 93.570 3.670 99.170 4.280 ;
        RECT 100.010 3.670 105.610 4.280 ;
      LAYER met3 ;
        RECT 3.990 108.480 105.400 108.965 ;
        RECT 3.990 107.120 105.000 108.480 ;
        RECT 4.400 107.080 105.000 107.120 ;
        RECT 4.400 105.720 105.400 107.080 ;
        RECT 3.990 100.320 105.400 105.720 ;
        RECT 3.990 98.920 105.000 100.320 ;
        RECT 3.990 92.160 105.400 98.920 ;
        RECT 3.990 90.760 105.000 92.160 ;
        RECT 3.990 88.080 105.400 90.760 ;
        RECT 4.400 86.680 105.400 88.080 ;
        RECT 3.990 84.000 105.400 86.680 ;
        RECT 3.990 82.600 105.000 84.000 ;
        RECT 3.990 75.840 105.400 82.600 ;
        RECT 3.990 74.440 105.000 75.840 ;
        RECT 3.990 69.040 105.400 74.440 ;
        RECT 4.400 67.680 105.400 69.040 ;
        RECT 4.400 67.640 105.000 67.680 ;
        RECT 3.990 66.280 105.000 67.640 ;
        RECT 3.990 59.520 105.400 66.280 ;
        RECT 3.990 58.120 105.000 59.520 ;
        RECT 3.990 51.360 105.400 58.120 ;
        RECT 3.990 50.000 105.000 51.360 ;
        RECT 4.400 49.960 105.000 50.000 ;
        RECT 4.400 48.600 105.400 49.960 ;
        RECT 3.990 43.200 105.400 48.600 ;
        RECT 3.990 41.800 105.000 43.200 ;
        RECT 3.990 35.040 105.400 41.800 ;
        RECT 3.990 33.640 105.000 35.040 ;
        RECT 3.990 30.960 105.400 33.640 ;
        RECT 4.400 29.560 105.400 30.960 ;
        RECT 3.990 26.880 105.400 29.560 ;
        RECT 3.990 25.480 105.000 26.880 ;
        RECT 3.990 18.720 105.400 25.480 ;
        RECT 3.990 17.320 105.000 18.720 ;
        RECT 3.990 11.920 105.400 17.320 ;
        RECT 4.400 10.560 105.400 11.920 ;
        RECT 4.400 10.520 105.000 10.560 ;
        RECT 3.990 9.695 105.000 10.520 ;
  END
END digital
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1754794521
<< error_p >>
rect -653 246 -595 252
rect -461 246 -403 252
rect -269 246 -211 252
rect -77 246 -19 252
rect 115 246 173 252
rect 307 246 365 252
rect 499 246 557 252
rect 691 246 749 252
rect -653 212 -641 246
rect -461 212 -449 246
rect -269 212 -257 246
rect -77 212 -65 246
rect 115 212 127 246
rect 307 212 319 246
rect 499 212 511 246
rect 691 212 703 246
rect -653 206 -595 212
rect -461 206 -403 212
rect -269 206 -211 212
rect -77 206 -19 212
rect 115 206 173 212
rect 307 206 365 212
rect 499 206 557 212
rect 691 206 749 212
rect -749 -212 -691 -206
rect -557 -212 -499 -206
rect -365 -212 -307 -206
rect -173 -212 -115 -206
rect 19 -212 77 -206
rect 211 -212 269 -206
rect 403 -212 461 -206
rect 595 -212 653 -206
rect -749 -246 -737 -212
rect -557 -246 -545 -212
rect -365 -246 -353 -212
rect -173 -246 -161 -212
rect 19 -246 31 -212
rect 211 -246 223 -212
rect 403 -246 415 -212
rect 595 -246 607 -212
rect -749 -252 -691 -246
rect -557 -252 -499 -246
rect -365 -252 -307 -246
rect -173 -252 -115 -246
rect 19 -252 77 -246
rect 211 -252 269 -246
rect 403 -252 461 -246
rect 595 -252 653 -246
<< nwell >>
rect -737 227 833 265
rect -833 -227 833 227
rect -833 -265 737 -227
<< pmos >>
rect -735 -165 -705 165
rect -639 -165 -609 165
rect -543 -165 -513 165
rect -447 -165 -417 165
rect -351 -165 -321 165
rect -255 -165 -225 165
rect -159 -165 -129 165
rect -63 -165 -33 165
rect 33 -165 63 165
rect 129 -165 159 165
rect 225 -165 255 165
rect 321 -165 351 165
rect 417 -165 447 165
rect 513 -165 543 165
rect 609 -165 639 165
rect 705 -165 735 165
<< pdiff >>
rect -797 153 -735 165
rect -797 -153 -785 153
rect -751 -153 -735 153
rect -797 -165 -735 -153
rect -705 153 -639 165
rect -705 -153 -689 153
rect -655 -153 -639 153
rect -705 -165 -639 -153
rect -609 153 -543 165
rect -609 -153 -593 153
rect -559 -153 -543 153
rect -609 -165 -543 -153
rect -513 153 -447 165
rect -513 -153 -497 153
rect -463 -153 -447 153
rect -513 -165 -447 -153
rect -417 153 -351 165
rect -417 -153 -401 153
rect -367 -153 -351 153
rect -417 -165 -351 -153
rect -321 153 -255 165
rect -321 -153 -305 153
rect -271 -153 -255 153
rect -321 -165 -255 -153
rect -225 153 -159 165
rect -225 -153 -209 153
rect -175 -153 -159 153
rect -225 -165 -159 -153
rect -129 153 -63 165
rect -129 -153 -113 153
rect -79 -153 -63 153
rect -129 -165 -63 -153
rect -33 153 33 165
rect -33 -153 -17 153
rect 17 -153 33 153
rect -33 -165 33 -153
rect 63 153 129 165
rect 63 -153 79 153
rect 113 -153 129 153
rect 63 -165 129 -153
rect 159 153 225 165
rect 159 -153 175 153
rect 209 -153 225 153
rect 159 -165 225 -153
rect 255 153 321 165
rect 255 -153 271 153
rect 305 -153 321 153
rect 255 -165 321 -153
rect 351 153 417 165
rect 351 -153 367 153
rect 401 -153 417 153
rect 351 -165 417 -153
rect 447 153 513 165
rect 447 -153 463 153
rect 497 -153 513 153
rect 447 -165 513 -153
rect 543 153 609 165
rect 543 -153 559 153
rect 593 -153 609 153
rect 543 -165 609 -153
rect 639 153 705 165
rect 639 -153 655 153
rect 689 -153 705 153
rect 639 -165 705 -153
rect 735 153 797 165
rect 735 -153 751 153
rect 785 -153 797 153
rect 735 -165 797 -153
<< pdiffc >>
rect -785 -153 -751 153
rect -689 -153 -655 153
rect -593 -153 -559 153
rect -497 -153 -463 153
rect -401 -153 -367 153
rect -305 -153 -271 153
rect -209 -153 -175 153
rect -113 -153 -79 153
rect -17 -153 17 153
rect 79 -153 113 153
rect 175 -153 209 153
rect 271 -153 305 153
rect 367 -153 401 153
rect 463 -153 497 153
rect 559 -153 593 153
rect 655 -153 689 153
rect 751 -153 785 153
<< poly >>
rect -657 246 -591 262
rect -657 212 -641 246
rect -607 212 -591 246
rect -657 196 -591 212
rect -465 246 -399 262
rect -465 212 -449 246
rect -415 212 -399 246
rect -465 196 -399 212
rect -273 246 -207 262
rect -273 212 -257 246
rect -223 212 -207 246
rect -273 196 -207 212
rect -81 246 -15 262
rect -81 212 -65 246
rect -31 212 -15 246
rect -81 196 -15 212
rect 111 246 177 262
rect 111 212 127 246
rect 161 212 177 246
rect 111 196 177 212
rect 303 246 369 262
rect 303 212 319 246
rect 353 212 369 246
rect 303 196 369 212
rect 495 246 561 262
rect 495 212 511 246
rect 545 212 561 246
rect 495 196 561 212
rect 687 246 753 262
rect 687 212 703 246
rect 737 212 753 246
rect 687 196 753 212
rect -735 165 -705 191
rect -639 165 -609 196
rect -543 165 -513 191
rect -447 165 -417 196
rect -351 165 -321 191
rect -255 165 -225 196
rect -159 165 -129 191
rect -63 165 -33 196
rect 33 165 63 191
rect 129 165 159 196
rect 225 165 255 191
rect 321 165 351 196
rect 417 165 447 191
rect 513 165 543 196
rect 609 165 639 191
rect 705 165 735 196
rect -735 -196 -705 -165
rect -639 -191 -609 -165
rect -543 -196 -513 -165
rect -447 -191 -417 -165
rect -351 -196 -321 -165
rect -255 -191 -225 -165
rect -159 -196 -129 -165
rect -63 -191 -33 -165
rect 33 -196 63 -165
rect 129 -191 159 -165
rect 225 -196 255 -165
rect 321 -191 351 -165
rect 417 -196 447 -165
rect 513 -191 543 -165
rect 609 -196 639 -165
rect 705 -191 735 -165
rect -753 -212 -687 -196
rect -753 -246 -737 -212
rect -703 -246 -687 -212
rect -753 -262 -687 -246
rect -561 -212 -495 -196
rect -561 -246 -545 -212
rect -511 -246 -495 -212
rect -561 -262 -495 -246
rect -369 -212 -303 -196
rect -369 -246 -353 -212
rect -319 -246 -303 -212
rect -369 -262 -303 -246
rect -177 -212 -111 -196
rect -177 -246 -161 -212
rect -127 -246 -111 -212
rect -177 -262 -111 -246
rect 15 -212 81 -196
rect 15 -246 31 -212
rect 65 -246 81 -212
rect 15 -262 81 -246
rect 207 -212 273 -196
rect 207 -246 223 -212
rect 257 -246 273 -212
rect 207 -262 273 -246
rect 399 -212 465 -196
rect 399 -246 415 -212
rect 449 -246 465 -212
rect 399 -262 465 -246
rect 591 -212 657 -196
rect 591 -246 607 -212
rect 641 -246 657 -212
rect 591 -262 657 -246
<< polycont >>
rect -641 212 -607 246
rect -449 212 -415 246
rect -257 212 -223 246
rect -65 212 -31 246
rect 127 212 161 246
rect 319 212 353 246
rect 511 212 545 246
rect 703 212 737 246
rect -737 -246 -703 -212
rect -545 -246 -511 -212
rect -353 -246 -319 -212
rect -161 -246 -127 -212
rect 31 -246 65 -212
rect 223 -246 257 -212
rect 415 -246 449 -212
rect 607 -246 641 -212
<< locali >>
rect -657 212 -641 246
rect -607 212 -591 246
rect -465 212 -449 246
rect -415 212 -399 246
rect -273 212 -257 246
rect -223 212 -207 246
rect -81 212 -65 246
rect -31 212 -15 246
rect 111 212 127 246
rect 161 212 177 246
rect 303 212 319 246
rect 353 212 369 246
rect 495 212 511 246
rect 545 212 561 246
rect 687 212 703 246
rect 737 212 753 246
rect -785 153 -751 169
rect -785 -169 -751 -153
rect -689 153 -655 169
rect -689 -169 -655 -153
rect -593 153 -559 169
rect -593 -169 -559 -153
rect -497 153 -463 169
rect -497 -169 -463 -153
rect -401 153 -367 169
rect -401 -169 -367 -153
rect -305 153 -271 169
rect -305 -169 -271 -153
rect -209 153 -175 169
rect -209 -169 -175 -153
rect -113 153 -79 169
rect -113 -169 -79 -153
rect -17 153 17 169
rect -17 -169 17 -153
rect 79 153 113 169
rect 79 -169 113 -153
rect 175 153 209 169
rect 175 -169 209 -153
rect 271 153 305 169
rect 271 -169 305 -153
rect 367 153 401 169
rect 367 -169 401 -153
rect 463 153 497 169
rect 463 -169 497 -153
rect 559 153 593 169
rect 559 -169 593 -153
rect 655 153 689 169
rect 655 -169 689 -153
rect 751 153 785 169
rect 751 -169 785 -153
rect -753 -246 -737 -212
rect -703 -246 -687 -212
rect -561 -246 -545 -212
rect -511 -246 -495 -212
rect -369 -246 -353 -212
rect -319 -246 -303 -212
rect -177 -246 -161 -212
rect -127 -246 -111 -212
rect 15 -246 31 -212
rect 65 -246 81 -212
rect 207 -246 223 -212
rect 257 -246 273 -212
rect 399 -246 415 -212
rect 449 -246 465 -212
rect 591 -246 607 -212
rect 641 -246 657 -212
<< viali >>
rect -641 212 -607 246
rect -449 212 -415 246
rect -257 212 -223 246
rect -65 212 -31 246
rect 127 212 161 246
rect 319 212 353 246
rect 511 212 545 246
rect 703 212 737 246
rect -785 44 -751 136
rect -689 -136 -655 -44
rect -593 44 -559 136
rect -497 -136 -463 -44
rect -401 44 -367 136
rect -305 -136 -271 -44
rect -209 44 -175 136
rect -113 -136 -79 -44
rect -17 44 17 136
rect 79 -136 113 -44
rect 175 44 209 136
rect 271 -136 305 -44
rect 367 44 401 136
rect 463 -136 497 -44
rect 559 44 593 136
rect 655 -136 689 -44
rect 751 44 785 136
rect -737 -246 -703 -212
rect -545 -246 -511 -212
rect -353 -246 -319 -212
rect -161 -246 -127 -212
rect 31 -246 65 -212
rect 223 -246 257 -212
rect 415 -246 449 -212
rect 607 -246 641 -212
<< metal1 >>
rect -653 246 -595 252
rect -653 212 -641 246
rect -607 212 -595 246
rect -653 206 -595 212
rect -461 246 -403 252
rect -461 212 -449 246
rect -415 212 -403 246
rect -461 206 -403 212
rect -269 246 -211 252
rect -269 212 -257 246
rect -223 212 -211 246
rect -269 206 -211 212
rect -77 246 -19 252
rect -77 212 -65 246
rect -31 212 -19 246
rect -77 206 -19 212
rect 115 246 173 252
rect 115 212 127 246
rect 161 212 173 246
rect 115 206 173 212
rect 307 246 365 252
rect 307 212 319 246
rect 353 212 365 246
rect 307 206 365 212
rect 499 246 557 252
rect 499 212 511 246
rect 545 212 557 246
rect 499 206 557 212
rect 691 246 749 252
rect 691 212 703 246
rect 737 212 749 246
rect 691 206 749 212
rect -791 136 -745 148
rect -791 44 -785 136
rect -751 44 -745 136
rect -791 32 -745 44
rect -599 136 -553 148
rect -599 44 -593 136
rect -559 44 -553 136
rect -599 32 -553 44
rect -407 136 -361 148
rect -407 44 -401 136
rect -367 44 -361 136
rect -407 32 -361 44
rect -215 136 -169 148
rect -215 44 -209 136
rect -175 44 -169 136
rect -215 32 -169 44
rect -23 136 23 148
rect -23 44 -17 136
rect 17 44 23 136
rect -23 32 23 44
rect 169 136 215 148
rect 169 44 175 136
rect 209 44 215 136
rect 169 32 215 44
rect 361 136 407 148
rect 361 44 367 136
rect 401 44 407 136
rect 361 32 407 44
rect 553 136 599 148
rect 553 44 559 136
rect 593 44 599 136
rect 553 32 599 44
rect 745 136 791 148
rect 745 44 751 136
rect 785 44 791 136
rect 745 32 791 44
rect -695 -44 -649 -32
rect -695 -136 -689 -44
rect -655 -136 -649 -44
rect -695 -148 -649 -136
rect -503 -44 -457 -32
rect -503 -136 -497 -44
rect -463 -136 -457 -44
rect -503 -148 -457 -136
rect -311 -44 -265 -32
rect -311 -136 -305 -44
rect -271 -136 -265 -44
rect -311 -148 -265 -136
rect -119 -44 -73 -32
rect -119 -136 -113 -44
rect -79 -136 -73 -44
rect -119 -148 -73 -136
rect 73 -44 119 -32
rect 73 -136 79 -44
rect 113 -136 119 -44
rect 73 -148 119 -136
rect 265 -44 311 -32
rect 265 -136 271 -44
rect 305 -136 311 -44
rect 265 -148 311 -136
rect 457 -44 503 -32
rect 457 -136 463 -44
rect 497 -136 503 -44
rect 457 -148 503 -136
rect 649 -44 695 -32
rect 649 -136 655 -44
rect 689 -136 695 -44
rect 649 -148 695 -136
rect -749 -212 -691 -206
rect -749 -246 -737 -212
rect -703 -246 -691 -212
rect -749 -252 -691 -246
rect -557 -212 -499 -206
rect -557 -246 -545 -212
rect -511 -246 -499 -212
rect -557 -252 -499 -246
rect -365 -212 -307 -206
rect -365 -246 -353 -212
rect -319 -246 -307 -212
rect -365 -252 -307 -246
rect -173 -212 -115 -206
rect -173 -246 -161 -212
rect -127 -246 -115 -212
rect -173 -252 -115 -246
rect 19 -212 77 -206
rect 19 -246 31 -212
rect 65 -246 77 -212
rect 19 -252 77 -246
rect 211 -212 269 -206
rect 211 -246 223 -212
rect 257 -246 269 -212
rect 211 -252 269 -246
rect 403 -212 461 -206
rect 403 -246 415 -212
rect 449 -246 461 -212
rect 403 -252 461 -246
rect 595 -212 653 -206
rect 595 -246 607 -212
rect 641 -246 653 -212
rect 595 -252 653 -246
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.65 l 0.15 m 1 nf 16 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc +30 viadrn -30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1755037679
<< metal3 >>
rect -3104 5132 -1732 5160
rect -3104 4108 -1816 5132
rect -1752 4108 -1732 5132
rect -3104 4080 -1732 4108
rect -1492 5132 -120 5160
rect -1492 4108 -204 5132
rect -140 4108 -120 5132
rect -1492 4080 -120 4108
rect 120 5132 1492 5160
rect 120 4108 1408 5132
rect 1472 4108 1492 5132
rect 120 4080 1492 4108
rect 1732 5132 3104 5160
rect 1732 4108 3020 5132
rect 3084 4108 3104 5132
rect 1732 4080 3104 4108
rect -3104 3812 -1732 3840
rect -3104 2788 -1816 3812
rect -1752 2788 -1732 3812
rect -3104 2760 -1732 2788
rect -1492 3812 -120 3840
rect -1492 2788 -204 3812
rect -140 2788 -120 3812
rect -1492 2760 -120 2788
rect 120 3812 1492 3840
rect 120 2788 1408 3812
rect 1472 2788 1492 3812
rect 120 2760 1492 2788
rect 1732 3812 3104 3840
rect 1732 2788 3020 3812
rect 3084 2788 3104 3812
rect 1732 2760 3104 2788
rect -3104 2492 -1732 2520
rect -3104 1468 -1816 2492
rect -1752 1468 -1732 2492
rect -3104 1440 -1732 1468
rect -1492 2492 -120 2520
rect -1492 1468 -204 2492
rect -140 1468 -120 2492
rect -1492 1440 -120 1468
rect 120 2492 1492 2520
rect 120 1468 1408 2492
rect 1472 1468 1492 2492
rect 120 1440 1492 1468
rect 1732 2492 3104 2520
rect 1732 1468 3020 2492
rect 3084 1468 3104 2492
rect 1732 1440 3104 1468
rect -3104 1172 -1732 1200
rect -3104 148 -1816 1172
rect -1752 148 -1732 1172
rect -3104 120 -1732 148
rect -1492 1172 -120 1200
rect -1492 148 -204 1172
rect -140 148 -120 1172
rect -1492 120 -120 148
rect 120 1172 1492 1200
rect 120 148 1408 1172
rect 1472 148 1492 1172
rect 120 120 1492 148
rect 1732 1172 3104 1200
rect 1732 148 3020 1172
rect 3084 148 3104 1172
rect 1732 120 3104 148
rect -3104 -148 -1732 -120
rect -3104 -1172 -1816 -148
rect -1752 -1172 -1732 -148
rect -3104 -1200 -1732 -1172
rect -1492 -148 -120 -120
rect -1492 -1172 -204 -148
rect -140 -1172 -120 -148
rect -1492 -1200 -120 -1172
rect 120 -148 1492 -120
rect 120 -1172 1408 -148
rect 1472 -1172 1492 -148
rect 120 -1200 1492 -1172
rect 1732 -148 3104 -120
rect 1732 -1172 3020 -148
rect 3084 -1172 3104 -148
rect 1732 -1200 3104 -1172
rect -3104 -1468 -1732 -1440
rect -3104 -2492 -1816 -1468
rect -1752 -2492 -1732 -1468
rect -3104 -2520 -1732 -2492
rect -1492 -1468 -120 -1440
rect -1492 -2492 -204 -1468
rect -140 -2492 -120 -1468
rect -1492 -2520 -120 -2492
rect 120 -1468 1492 -1440
rect 120 -2492 1408 -1468
rect 1472 -2492 1492 -1468
rect 120 -2520 1492 -2492
rect 1732 -1468 3104 -1440
rect 1732 -2492 3020 -1468
rect 3084 -2492 3104 -1468
rect 1732 -2520 3104 -2492
rect -3104 -2788 -1732 -2760
rect -3104 -3812 -1816 -2788
rect -1752 -3812 -1732 -2788
rect -3104 -3840 -1732 -3812
rect -1492 -2788 -120 -2760
rect -1492 -3812 -204 -2788
rect -140 -3812 -120 -2788
rect -1492 -3840 -120 -3812
rect 120 -2788 1492 -2760
rect 120 -3812 1408 -2788
rect 1472 -3812 1492 -2788
rect 120 -3840 1492 -3812
rect 1732 -2788 3104 -2760
rect 1732 -3812 3020 -2788
rect 3084 -3812 3104 -2788
rect 1732 -3840 3104 -3812
rect -3104 -4108 -1732 -4080
rect -3104 -5132 -1816 -4108
rect -1752 -5132 -1732 -4108
rect -3104 -5160 -1732 -5132
rect -1492 -4108 -120 -4080
rect -1492 -5132 -204 -4108
rect -140 -5132 -120 -4108
rect -1492 -5160 -120 -5132
rect 120 -4108 1492 -4080
rect 120 -5132 1408 -4108
rect 1472 -5132 1492 -4108
rect 120 -5160 1492 -5132
rect 1732 -4108 3104 -4080
rect 1732 -5132 3020 -4108
rect 3084 -5132 3104 -4108
rect 1732 -5160 3104 -5132
<< via3 >>
rect -1816 4108 -1752 5132
rect -204 4108 -140 5132
rect 1408 4108 1472 5132
rect 3020 4108 3084 5132
rect -1816 2788 -1752 3812
rect -204 2788 -140 3812
rect 1408 2788 1472 3812
rect 3020 2788 3084 3812
rect -1816 1468 -1752 2492
rect -204 1468 -140 2492
rect 1408 1468 1472 2492
rect 3020 1468 3084 2492
rect -1816 148 -1752 1172
rect -204 148 -140 1172
rect 1408 148 1472 1172
rect 3020 148 3084 1172
rect -1816 -1172 -1752 -148
rect -204 -1172 -140 -148
rect 1408 -1172 1472 -148
rect 3020 -1172 3084 -148
rect -1816 -2492 -1752 -1468
rect -204 -2492 -140 -1468
rect 1408 -2492 1472 -1468
rect 3020 -2492 3084 -1468
rect -1816 -3812 -1752 -2788
rect -204 -3812 -140 -2788
rect 1408 -3812 1472 -2788
rect 3020 -3812 3084 -2788
rect -1816 -5132 -1752 -4108
rect -204 -5132 -140 -4108
rect 1408 -5132 1472 -4108
rect 3020 -5132 3084 -4108
<< mimcap >>
rect -3064 5080 -2064 5120
rect -3064 4160 -3024 5080
rect -2104 4160 -2064 5080
rect -3064 4120 -2064 4160
rect -1452 5080 -452 5120
rect -1452 4160 -1412 5080
rect -492 4160 -452 5080
rect -1452 4120 -452 4160
rect 160 5080 1160 5120
rect 160 4160 200 5080
rect 1120 4160 1160 5080
rect 160 4120 1160 4160
rect 1772 5080 2772 5120
rect 1772 4160 1812 5080
rect 2732 4160 2772 5080
rect 1772 4120 2772 4160
rect -3064 3760 -2064 3800
rect -3064 2840 -3024 3760
rect -2104 2840 -2064 3760
rect -3064 2800 -2064 2840
rect -1452 3760 -452 3800
rect -1452 2840 -1412 3760
rect -492 2840 -452 3760
rect -1452 2800 -452 2840
rect 160 3760 1160 3800
rect 160 2840 200 3760
rect 1120 2840 1160 3760
rect 160 2800 1160 2840
rect 1772 3760 2772 3800
rect 1772 2840 1812 3760
rect 2732 2840 2772 3760
rect 1772 2800 2772 2840
rect -3064 2440 -2064 2480
rect -3064 1520 -3024 2440
rect -2104 1520 -2064 2440
rect -3064 1480 -2064 1520
rect -1452 2440 -452 2480
rect -1452 1520 -1412 2440
rect -492 1520 -452 2440
rect -1452 1480 -452 1520
rect 160 2440 1160 2480
rect 160 1520 200 2440
rect 1120 1520 1160 2440
rect 160 1480 1160 1520
rect 1772 2440 2772 2480
rect 1772 1520 1812 2440
rect 2732 1520 2772 2440
rect 1772 1480 2772 1520
rect -3064 1120 -2064 1160
rect -3064 200 -3024 1120
rect -2104 200 -2064 1120
rect -3064 160 -2064 200
rect -1452 1120 -452 1160
rect -1452 200 -1412 1120
rect -492 200 -452 1120
rect -1452 160 -452 200
rect 160 1120 1160 1160
rect 160 200 200 1120
rect 1120 200 1160 1120
rect 160 160 1160 200
rect 1772 1120 2772 1160
rect 1772 200 1812 1120
rect 2732 200 2772 1120
rect 1772 160 2772 200
rect -3064 -200 -2064 -160
rect -3064 -1120 -3024 -200
rect -2104 -1120 -2064 -200
rect -3064 -1160 -2064 -1120
rect -1452 -200 -452 -160
rect -1452 -1120 -1412 -200
rect -492 -1120 -452 -200
rect -1452 -1160 -452 -1120
rect 160 -200 1160 -160
rect 160 -1120 200 -200
rect 1120 -1120 1160 -200
rect 160 -1160 1160 -1120
rect 1772 -200 2772 -160
rect 1772 -1120 1812 -200
rect 2732 -1120 2772 -200
rect 1772 -1160 2772 -1120
rect -3064 -1520 -2064 -1480
rect -3064 -2440 -3024 -1520
rect -2104 -2440 -2064 -1520
rect -3064 -2480 -2064 -2440
rect -1452 -1520 -452 -1480
rect -1452 -2440 -1412 -1520
rect -492 -2440 -452 -1520
rect -1452 -2480 -452 -2440
rect 160 -1520 1160 -1480
rect 160 -2440 200 -1520
rect 1120 -2440 1160 -1520
rect 160 -2480 1160 -2440
rect 1772 -1520 2772 -1480
rect 1772 -2440 1812 -1520
rect 2732 -2440 2772 -1520
rect 1772 -2480 2772 -2440
rect -3064 -2840 -2064 -2800
rect -3064 -3760 -3024 -2840
rect -2104 -3760 -2064 -2840
rect -3064 -3800 -2064 -3760
rect -1452 -2840 -452 -2800
rect -1452 -3760 -1412 -2840
rect -492 -3760 -452 -2840
rect -1452 -3800 -452 -3760
rect 160 -2840 1160 -2800
rect 160 -3760 200 -2840
rect 1120 -3760 1160 -2840
rect 160 -3800 1160 -3760
rect 1772 -2840 2772 -2800
rect 1772 -3760 1812 -2840
rect 2732 -3760 2772 -2840
rect 1772 -3800 2772 -3760
rect -3064 -4160 -2064 -4120
rect -3064 -5080 -3024 -4160
rect -2104 -5080 -2064 -4160
rect -3064 -5120 -2064 -5080
rect -1452 -4160 -452 -4120
rect -1452 -5080 -1412 -4160
rect -492 -5080 -452 -4160
rect -1452 -5120 -452 -5080
rect 160 -4160 1160 -4120
rect 160 -5080 200 -4160
rect 1120 -5080 1160 -4160
rect 160 -5120 1160 -5080
rect 1772 -4160 2772 -4120
rect 1772 -5080 1812 -4160
rect 2732 -5080 2772 -4160
rect 1772 -5120 2772 -5080
<< mimcapcontact >>
rect -3024 4160 -2104 5080
rect -1412 4160 -492 5080
rect 200 4160 1120 5080
rect 1812 4160 2732 5080
rect -3024 2840 -2104 3760
rect -1412 2840 -492 3760
rect 200 2840 1120 3760
rect 1812 2840 2732 3760
rect -3024 1520 -2104 2440
rect -1412 1520 -492 2440
rect 200 1520 1120 2440
rect 1812 1520 2732 2440
rect -3024 200 -2104 1120
rect -1412 200 -492 1120
rect 200 200 1120 1120
rect 1812 200 2732 1120
rect -3024 -1120 -2104 -200
rect -1412 -1120 -492 -200
rect 200 -1120 1120 -200
rect 1812 -1120 2732 -200
rect -3024 -2440 -2104 -1520
rect -1412 -2440 -492 -1520
rect 200 -2440 1120 -1520
rect 1812 -2440 2732 -1520
rect -3024 -3760 -2104 -2840
rect -1412 -3760 -492 -2840
rect 200 -3760 1120 -2840
rect 1812 -3760 2732 -2840
rect -3024 -5080 -2104 -4160
rect -1412 -5080 -492 -4160
rect 200 -5080 1120 -4160
rect 1812 -5080 2732 -4160
<< metal4 >>
rect -2616 5081 -2512 5280
rect -1836 5132 -1732 5280
rect -3025 5080 -2103 5081
rect -3025 4160 -3024 5080
rect -2104 4160 -2103 5080
rect -3025 4159 -2103 4160
rect -2616 3761 -2512 4159
rect -1836 4108 -1816 5132
rect -1752 4108 -1732 5132
rect -1004 5081 -900 5280
rect -224 5132 -120 5280
rect -1413 5080 -491 5081
rect -1413 4160 -1412 5080
rect -492 4160 -491 5080
rect -1413 4159 -491 4160
rect -1836 3812 -1732 4108
rect -3025 3760 -2103 3761
rect -3025 2840 -3024 3760
rect -2104 2840 -2103 3760
rect -3025 2839 -2103 2840
rect -2616 2441 -2512 2839
rect -1836 2788 -1816 3812
rect -1752 2788 -1732 3812
rect -1004 3761 -900 4159
rect -224 4108 -204 5132
rect -140 4108 -120 5132
rect 608 5081 712 5280
rect 1388 5132 1492 5280
rect 199 5080 1121 5081
rect 199 4160 200 5080
rect 1120 4160 1121 5080
rect 199 4159 1121 4160
rect -224 3812 -120 4108
rect -1413 3760 -491 3761
rect -1413 2840 -1412 3760
rect -492 2840 -491 3760
rect -1413 2839 -491 2840
rect -1836 2492 -1732 2788
rect -3025 2440 -2103 2441
rect -3025 1520 -3024 2440
rect -2104 1520 -2103 2440
rect -3025 1519 -2103 1520
rect -2616 1121 -2512 1519
rect -1836 1468 -1816 2492
rect -1752 1468 -1732 2492
rect -1004 2441 -900 2839
rect -224 2788 -204 3812
rect -140 2788 -120 3812
rect 608 3761 712 4159
rect 1388 4108 1408 5132
rect 1472 4108 1492 5132
rect 2220 5081 2324 5280
rect 3000 5132 3104 5280
rect 1811 5080 2733 5081
rect 1811 4160 1812 5080
rect 2732 4160 2733 5080
rect 1811 4159 2733 4160
rect 1388 3812 1492 4108
rect 199 3760 1121 3761
rect 199 2840 200 3760
rect 1120 2840 1121 3760
rect 199 2839 1121 2840
rect -224 2492 -120 2788
rect -1413 2440 -491 2441
rect -1413 1520 -1412 2440
rect -492 1520 -491 2440
rect -1413 1519 -491 1520
rect -1836 1172 -1732 1468
rect -3025 1120 -2103 1121
rect -3025 200 -3024 1120
rect -2104 200 -2103 1120
rect -3025 199 -2103 200
rect -2616 -199 -2512 199
rect -1836 148 -1816 1172
rect -1752 148 -1732 1172
rect -1004 1121 -900 1519
rect -224 1468 -204 2492
rect -140 1468 -120 2492
rect 608 2441 712 2839
rect 1388 2788 1408 3812
rect 1472 2788 1492 3812
rect 2220 3761 2324 4159
rect 3000 4108 3020 5132
rect 3084 4108 3104 5132
rect 3000 3812 3104 4108
rect 1811 3760 2733 3761
rect 1811 2840 1812 3760
rect 2732 2840 2733 3760
rect 1811 2839 2733 2840
rect 1388 2492 1492 2788
rect 199 2440 1121 2441
rect 199 1520 200 2440
rect 1120 1520 1121 2440
rect 199 1519 1121 1520
rect -224 1172 -120 1468
rect -1413 1120 -491 1121
rect -1413 200 -1412 1120
rect -492 200 -491 1120
rect -1413 199 -491 200
rect -1836 -148 -1732 148
rect -3025 -200 -2103 -199
rect -3025 -1120 -3024 -200
rect -2104 -1120 -2103 -200
rect -3025 -1121 -2103 -1120
rect -2616 -1519 -2512 -1121
rect -1836 -1172 -1816 -148
rect -1752 -1172 -1732 -148
rect -1004 -199 -900 199
rect -224 148 -204 1172
rect -140 148 -120 1172
rect 608 1121 712 1519
rect 1388 1468 1408 2492
rect 1472 1468 1492 2492
rect 2220 2441 2324 2839
rect 3000 2788 3020 3812
rect 3084 2788 3104 3812
rect 3000 2492 3104 2788
rect 1811 2440 2733 2441
rect 1811 1520 1812 2440
rect 2732 1520 2733 2440
rect 1811 1519 2733 1520
rect 1388 1172 1492 1468
rect 199 1120 1121 1121
rect 199 200 200 1120
rect 1120 200 1121 1120
rect 199 199 1121 200
rect -224 -148 -120 148
rect -1413 -200 -491 -199
rect -1413 -1120 -1412 -200
rect -492 -1120 -491 -200
rect -1413 -1121 -491 -1120
rect -1836 -1468 -1732 -1172
rect -3025 -1520 -2103 -1519
rect -3025 -2440 -3024 -1520
rect -2104 -2440 -2103 -1520
rect -3025 -2441 -2103 -2440
rect -2616 -2839 -2512 -2441
rect -1836 -2492 -1816 -1468
rect -1752 -2492 -1732 -1468
rect -1004 -1519 -900 -1121
rect -224 -1172 -204 -148
rect -140 -1172 -120 -148
rect 608 -199 712 199
rect 1388 148 1408 1172
rect 1472 148 1492 1172
rect 2220 1121 2324 1519
rect 3000 1468 3020 2492
rect 3084 1468 3104 2492
rect 3000 1172 3104 1468
rect 1811 1120 2733 1121
rect 1811 200 1812 1120
rect 2732 200 2733 1120
rect 1811 199 2733 200
rect 1388 -148 1492 148
rect 199 -200 1121 -199
rect 199 -1120 200 -200
rect 1120 -1120 1121 -200
rect 199 -1121 1121 -1120
rect -224 -1468 -120 -1172
rect -1413 -1520 -491 -1519
rect -1413 -2440 -1412 -1520
rect -492 -2440 -491 -1520
rect -1413 -2441 -491 -2440
rect -1836 -2788 -1732 -2492
rect -3025 -2840 -2103 -2839
rect -3025 -3760 -3024 -2840
rect -2104 -3760 -2103 -2840
rect -3025 -3761 -2103 -3760
rect -2616 -4159 -2512 -3761
rect -1836 -3812 -1816 -2788
rect -1752 -3812 -1732 -2788
rect -1004 -2839 -900 -2441
rect -224 -2492 -204 -1468
rect -140 -2492 -120 -1468
rect 608 -1519 712 -1121
rect 1388 -1172 1408 -148
rect 1472 -1172 1492 -148
rect 2220 -199 2324 199
rect 3000 148 3020 1172
rect 3084 148 3104 1172
rect 3000 -148 3104 148
rect 1811 -200 2733 -199
rect 1811 -1120 1812 -200
rect 2732 -1120 2733 -200
rect 1811 -1121 2733 -1120
rect 1388 -1468 1492 -1172
rect 199 -1520 1121 -1519
rect 199 -2440 200 -1520
rect 1120 -2440 1121 -1520
rect 199 -2441 1121 -2440
rect -224 -2788 -120 -2492
rect -1413 -2840 -491 -2839
rect -1413 -3760 -1412 -2840
rect -492 -3760 -491 -2840
rect -1413 -3761 -491 -3760
rect -1836 -4108 -1732 -3812
rect -3025 -4160 -2103 -4159
rect -3025 -5080 -3024 -4160
rect -2104 -5080 -2103 -4160
rect -3025 -5081 -2103 -5080
rect -2616 -5280 -2512 -5081
rect -1836 -5132 -1816 -4108
rect -1752 -5132 -1732 -4108
rect -1004 -4159 -900 -3761
rect -224 -3812 -204 -2788
rect -140 -3812 -120 -2788
rect 608 -2839 712 -2441
rect 1388 -2492 1408 -1468
rect 1472 -2492 1492 -1468
rect 2220 -1519 2324 -1121
rect 3000 -1172 3020 -148
rect 3084 -1172 3104 -148
rect 3000 -1468 3104 -1172
rect 1811 -1520 2733 -1519
rect 1811 -2440 1812 -1520
rect 2732 -2440 2733 -1520
rect 1811 -2441 2733 -2440
rect 1388 -2788 1492 -2492
rect 199 -2840 1121 -2839
rect 199 -3760 200 -2840
rect 1120 -3760 1121 -2840
rect 199 -3761 1121 -3760
rect -224 -4108 -120 -3812
rect -1413 -4160 -491 -4159
rect -1413 -5080 -1412 -4160
rect -492 -5080 -491 -4160
rect -1413 -5081 -491 -5080
rect -1836 -5280 -1732 -5132
rect -1004 -5280 -900 -5081
rect -224 -5132 -204 -4108
rect -140 -5132 -120 -4108
rect 608 -4159 712 -3761
rect 1388 -3812 1408 -2788
rect 1472 -3812 1492 -2788
rect 2220 -2839 2324 -2441
rect 3000 -2492 3020 -1468
rect 3084 -2492 3104 -1468
rect 3000 -2788 3104 -2492
rect 1811 -2840 2733 -2839
rect 1811 -3760 1812 -2840
rect 2732 -3760 2733 -2840
rect 1811 -3761 2733 -3760
rect 1388 -4108 1492 -3812
rect 199 -4160 1121 -4159
rect 199 -5080 200 -4160
rect 1120 -5080 1121 -4160
rect 199 -5081 1121 -5080
rect -224 -5280 -120 -5132
rect 608 -5280 712 -5081
rect 1388 -5132 1408 -4108
rect 1472 -5132 1492 -4108
rect 2220 -4159 2324 -3761
rect 3000 -3812 3020 -2788
rect 3084 -3812 3104 -2788
rect 3000 -4108 3104 -3812
rect 1811 -4160 2733 -4159
rect 1811 -5080 1812 -4160
rect 2732 -5080 2733 -4160
rect 1811 -5081 2733 -5080
rect 1388 -5280 1492 -5132
rect 2220 -5280 2324 -5081
rect 3000 -5132 3020 -4108
rect 3084 -5132 3104 -4108
rect 3000 -5280 3104 -5132
<< properties >>
string FIXED_BBOX 1732 4080 2812 5160
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5 l 5 val 53.8 carea 2.00 cperi 0.19 nx 4 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

magic
tech sky130A
timestamp 1754942031
<< end >>

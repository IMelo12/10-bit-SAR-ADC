magic
tech sky130A
magscale 1 2
timestamp 1754900058
<< metal3 >>
rect -12776 5132 -11404 5160
rect -12776 4108 -11488 5132
rect -11424 4108 -11404 5132
rect -12776 4080 -11404 4108
rect -11164 5132 -9792 5160
rect -11164 4108 -9876 5132
rect -9812 4108 -9792 5132
rect -11164 4080 -9792 4108
rect -9552 5132 -8180 5160
rect -9552 4108 -8264 5132
rect -8200 4108 -8180 5132
rect -9552 4080 -8180 4108
rect -7940 5132 -6568 5160
rect -7940 4108 -6652 5132
rect -6588 4108 -6568 5132
rect -7940 4080 -6568 4108
rect -6328 5132 -4956 5160
rect -6328 4108 -5040 5132
rect -4976 4108 -4956 5132
rect -6328 4080 -4956 4108
rect -4716 5132 -3344 5160
rect -4716 4108 -3428 5132
rect -3364 4108 -3344 5132
rect -4716 4080 -3344 4108
rect -3104 5132 -1732 5160
rect -3104 4108 -1816 5132
rect -1752 4108 -1732 5132
rect -3104 4080 -1732 4108
rect -1492 5132 -120 5160
rect -1492 4108 -204 5132
rect -140 4108 -120 5132
rect -1492 4080 -120 4108
rect 120 5132 1492 5160
rect 120 4108 1408 5132
rect 1472 4108 1492 5132
rect 120 4080 1492 4108
rect 1732 5132 3104 5160
rect 1732 4108 3020 5132
rect 3084 4108 3104 5132
rect 1732 4080 3104 4108
rect 3344 5132 4716 5160
rect 3344 4108 4632 5132
rect 4696 4108 4716 5132
rect 3344 4080 4716 4108
rect 4956 5132 6328 5160
rect 4956 4108 6244 5132
rect 6308 4108 6328 5132
rect 4956 4080 6328 4108
rect 6568 5132 7940 5160
rect 6568 4108 7856 5132
rect 7920 4108 7940 5132
rect 6568 4080 7940 4108
rect 8180 5132 9552 5160
rect 8180 4108 9468 5132
rect 9532 4108 9552 5132
rect 8180 4080 9552 4108
rect 9792 5132 11164 5160
rect 9792 4108 11080 5132
rect 11144 4108 11164 5132
rect 9792 4080 11164 4108
rect 11404 5132 12776 5160
rect 11404 4108 12692 5132
rect 12756 4108 12776 5132
rect 11404 4080 12776 4108
rect -12776 3812 -11404 3840
rect -12776 2788 -11488 3812
rect -11424 2788 -11404 3812
rect -12776 2760 -11404 2788
rect -11164 3812 -9792 3840
rect -11164 2788 -9876 3812
rect -9812 2788 -9792 3812
rect -11164 2760 -9792 2788
rect -9552 3812 -8180 3840
rect -9552 2788 -8264 3812
rect -8200 2788 -8180 3812
rect -9552 2760 -8180 2788
rect -7940 3812 -6568 3840
rect -7940 2788 -6652 3812
rect -6588 2788 -6568 3812
rect -7940 2760 -6568 2788
rect -6328 3812 -4956 3840
rect -6328 2788 -5040 3812
rect -4976 2788 -4956 3812
rect -6328 2760 -4956 2788
rect -4716 3812 -3344 3840
rect -4716 2788 -3428 3812
rect -3364 2788 -3344 3812
rect -4716 2760 -3344 2788
rect -3104 3812 -1732 3840
rect -3104 2788 -1816 3812
rect -1752 2788 -1732 3812
rect -3104 2760 -1732 2788
rect -1492 3812 -120 3840
rect -1492 2788 -204 3812
rect -140 2788 -120 3812
rect -1492 2760 -120 2788
rect 120 3812 1492 3840
rect 120 2788 1408 3812
rect 1472 2788 1492 3812
rect 120 2760 1492 2788
rect 1732 3812 3104 3840
rect 1732 2788 3020 3812
rect 3084 2788 3104 3812
rect 1732 2760 3104 2788
rect 3344 3812 4716 3840
rect 3344 2788 4632 3812
rect 4696 2788 4716 3812
rect 3344 2760 4716 2788
rect 4956 3812 6328 3840
rect 4956 2788 6244 3812
rect 6308 2788 6328 3812
rect 4956 2760 6328 2788
rect 6568 3812 7940 3840
rect 6568 2788 7856 3812
rect 7920 2788 7940 3812
rect 6568 2760 7940 2788
rect 8180 3812 9552 3840
rect 8180 2788 9468 3812
rect 9532 2788 9552 3812
rect 8180 2760 9552 2788
rect 9792 3812 11164 3840
rect 9792 2788 11080 3812
rect 11144 2788 11164 3812
rect 9792 2760 11164 2788
rect 11404 3812 12776 3840
rect 11404 2788 12692 3812
rect 12756 2788 12776 3812
rect 11404 2760 12776 2788
rect -12776 2492 -11404 2520
rect -12776 1468 -11488 2492
rect -11424 1468 -11404 2492
rect -12776 1440 -11404 1468
rect -11164 2492 -9792 2520
rect -11164 1468 -9876 2492
rect -9812 1468 -9792 2492
rect -11164 1440 -9792 1468
rect -9552 2492 -8180 2520
rect -9552 1468 -8264 2492
rect -8200 1468 -8180 2492
rect -9552 1440 -8180 1468
rect -7940 2492 -6568 2520
rect -7940 1468 -6652 2492
rect -6588 1468 -6568 2492
rect -7940 1440 -6568 1468
rect -6328 2492 -4956 2520
rect -6328 1468 -5040 2492
rect -4976 1468 -4956 2492
rect -6328 1440 -4956 1468
rect -4716 2492 -3344 2520
rect -4716 1468 -3428 2492
rect -3364 1468 -3344 2492
rect -4716 1440 -3344 1468
rect -3104 2492 -1732 2520
rect -3104 1468 -1816 2492
rect -1752 1468 -1732 2492
rect -3104 1440 -1732 1468
rect -1492 2492 -120 2520
rect -1492 1468 -204 2492
rect -140 1468 -120 2492
rect -1492 1440 -120 1468
rect 120 2492 1492 2520
rect 120 1468 1408 2492
rect 1472 1468 1492 2492
rect 120 1440 1492 1468
rect 1732 2492 3104 2520
rect 1732 1468 3020 2492
rect 3084 1468 3104 2492
rect 1732 1440 3104 1468
rect 3344 2492 4716 2520
rect 3344 1468 4632 2492
rect 4696 1468 4716 2492
rect 3344 1440 4716 1468
rect 4956 2492 6328 2520
rect 4956 1468 6244 2492
rect 6308 1468 6328 2492
rect 4956 1440 6328 1468
rect 6568 2492 7940 2520
rect 6568 1468 7856 2492
rect 7920 1468 7940 2492
rect 6568 1440 7940 1468
rect 8180 2492 9552 2520
rect 8180 1468 9468 2492
rect 9532 1468 9552 2492
rect 8180 1440 9552 1468
rect 9792 2492 11164 2520
rect 9792 1468 11080 2492
rect 11144 1468 11164 2492
rect 9792 1440 11164 1468
rect 11404 2492 12776 2520
rect 11404 1468 12692 2492
rect 12756 1468 12776 2492
rect 11404 1440 12776 1468
rect -12776 1172 -11404 1200
rect -12776 148 -11488 1172
rect -11424 148 -11404 1172
rect -12776 120 -11404 148
rect -11164 1172 -9792 1200
rect -11164 148 -9876 1172
rect -9812 148 -9792 1172
rect -11164 120 -9792 148
rect -9552 1172 -8180 1200
rect -9552 148 -8264 1172
rect -8200 148 -8180 1172
rect -9552 120 -8180 148
rect -7940 1172 -6568 1200
rect -7940 148 -6652 1172
rect -6588 148 -6568 1172
rect -7940 120 -6568 148
rect -6328 1172 -4956 1200
rect -6328 148 -5040 1172
rect -4976 148 -4956 1172
rect -6328 120 -4956 148
rect -4716 1172 -3344 1200
rect -4716 148 -3428 1172
rect -3364 148 -3344 1172
rect -4716 120 -3344 148
rect -3104 1172 -1732 1200
rect -3104 148 -1816 1172
rect -1752 148 -1732 1172
rect -3104 120 -1732 148
rect -1492 1172 -120 1200
rect -1492 148 -204 1172
rect -140 148 -120 1172
rect -1492 120 -120 148
rect 120 1172 1492 1200
rect 120 148 1408 1172
rect 1472 148 1492 1172
rect 120 120 1492 148
rect 1732 1172 3104 1200
rect 1732 148 3020 1172
rect 3084 148 3104 1172
rect 1732 120 3104 148
rect 3344 1172 4716 1200
rect 3344 148 4632 1172
rect 4696 148 4716 1172
rect 3344 120 4716 148
rect 4956 1172 6328 1200
rect 4956 148 6244 1172
rect 6308 148 6328 1172
rect 4956 120 6328 148
rect 6568 1172 7940 1200
rect 6568 148 7856 1172
rect 7920 148 7940 1172
rect 6568 120 7940 148
rect 8180 1172 9552 1200
rect 8180 148 9468 1172
rect 9532 148 9552 1172
rect 8180 120 9552 148
rect 9792 1172 11164 1200
rect 9792 148 11080 1172
rect 11144 148 11164 1172
rect 9792 120 11164 148
rect 11404 1172 12776 1200
rect 11404 148 12692 1172
rect 12756 148 12776 1172
rect 11404 120 12776 148
rect -12776 -148 -11404 -120
rect -12776 -1172 -11488 -148
rect -11424 -1172 -11404 -148
rect -12776 -1200 -11404 -1172
rect -11164 -148 -9792 -120
rect -11164 -1172 -9876 -148
rect -9812 -1172 -9792 -148
rect -11164 -1200 -9792 -1172
rect -9552 -148 -8180 -120
rect -9552 -1172 -8264 -148
rect -8200 -1172 -8180 -148
rect -9552 -1200 -8180 -1172
rect -7940 -148 -6568 -120
rect -7940 -1172 -6652 -148
rect -6588 -1172 -6568 -148
rect -7940 -1200 -6568 -1172
rect -6328 -148 -4956 -120
rect -6328 -1172 -5040 -148
rect -4976 -1172 -4956 -148
rect -6328 -1200 -4956 -1172
rect -4716 -148 -3344 -120
rect -4716 -1172 -3428 -148
rect -3364 -1172 -3344 -148
rect -4716 -1200 -3344 -1172
rect -3104 -148 -1732 -120
rect -3104 -1172 -1816 -148
rect -1752 -1172 -1732 -148
rect -3104 -1200 -1732 -1172
rect -1492 -148 -120 -120
rect -1492 -1172 -204 -148
rect -140 -1172 -120 -148
rect -1492 -1200 -120 -1172
rect 120 -148 1492 -120
rect 120 -1172 1408 -148
rect 1472 -1172 1492 -148
rect 120 -1200 1492 -1172
rect 1732 -148 3104 -120
rect 1732 -1172 3020 -148
rect 3084 -1172 3104 -148
rect 1732 -1200 3104 -1172
rect 3344 -148 4716 -120
rect 3344 -1172 4632 -148
rect 4696 -1172 4716 -148
rect 3344 -1200 4716 -1172
rect 4956 -148 6328 -120
rect 4956 -1172 6244 -148
rect 6308 -1172 6328 -148
rect 4956 -1200 6328 -1172
rect 6568 -148 7940 -120
rect 6568 -1172 7856 -148
rect 7920 -1172 7940 -148
rect 6568 -1200 7940 -1172
rect 8180 -148 9552 -120
rect 8180 -1172 9468 -148
rect 9532 -1172 9552 -148
rect 8180 -1200 9552 -1172
rect 9792 -148 11164 -120
rect 9792 -1172 11080 -148
rect 11144 -1172 11164 -148
rect 9792 -1200 11164 -1172
rect 11404 -148 12776 -120
rect 11404 -1172 12692 -148
rect 12756 -1172 12776 -148
rect 11404 -1200 12776 -1172
rect -12776 -1468 -11404 -1440
rect -12776 -2492 -11488 -1468
rect -11424 -2492 -11404 -1468
rect -12776 -2520 -11404 -2492
rect -11164 -1468 -9792 -1440
rect -11164 -2492 -9876 -1468
rect -9812 -2492 -9792 -1468
rect -11164 -2520 -9792 -2492
rect -9552 -1468 -8180 -1440
rect -9552 -2492 -8264 -1468
rect -8200 -2492 -8180 -1468
rect -9552 -2520 -8180 -2492
rect -7940 -1468 -6568 -1440
rect -7940 -2492 -6652 -1468
rect -6588 -2492 -6568 -1468
rect -7940 -2520 -6568 -2492
rect -6328 -1468 -4956 -1440
rect -6328 -2492 -5040 -1468
rect -4976 -2492 -4956 -1468
rect -6328 -2520 -4956 -2492
rect -4716 -1468 -3344 -1440
rect -4716 -2492 -3428 -1468
rect -3364 -2492 -3344 -1468
rect -4716 -2520 -3344 -2492
rect -3104 -1468 -1732 -1440
rect -3104 -2492 -1816 -1468
rect -1752 -2492 -1732 -1468
rect -3104 -2520 -1732 -2492
rect -1492 -1468 -120 -1440
rect -1492 -2492 -204 -1468
rect -140 -2492 -120 -1468
rect -1492 -2520 -120 -2492
rect 120 -1468 1492 -1440
rect 120 -2492 1408 -1468
rect 1472 -2492 1492 -1468
rect 120 -2520 1492 -2492
rect 1732 -1468 3104 -1440
rect 1732 -2492 3020 -1468
rect 3084 -2492 3104 -1468
rect 1732 -2520 3104 -2492
rect 3344 -1468 4716 -1440
rect 3344 -2492 4632 -1468
rect 4696 -2492 4716 -1468
rect 3344 -2520 4716 -2492
rect 4956 -1468 6328 -1440
rect 4956 -2492 6244 -1468
rect 6308 -2492 6328 -1468
rect 4956 -2520 6328 -2492
rect 6568 -1468 7940 -1440
rect 6568 -2492 7856 -1468
rect 7920 -2492 7940 -1468
rect 6568 -2520 7940 -2492
rect 8180 -1468 9552 -1440
rect 8180 -2492 9468 -1468
rect 9532 -2492 9552 -1468
rect 8180 -2520 9552 -2492
rect 9792 -1468 11164 -1440
rect 9792 -2492 11080 -1468
rect 11144 -2492 11164 -1468
rect 9792 -2520 11164 -2492
rect 11404 -1468 12776 -1440
rect 11404 -2492 12692 -1468
rect 12756 -2492 12776 -1468
rect 11404 -2520 12776 -2492
rect -12776 -2788 -11404 -2760
rect -12776 -3812 -11488 -2788
rect -11424 -3812 -11404 -2788
rect -12776 -3840 -11404 -3812
rect -11164 -2788 -9792 -2760
rect -11164 -3812 -9876 -2788
rect -9812 -3812 -9792 -2788
rect -11164 -3840 -9792 -3812
rect -9552 -2788 -8180 -2760
rect -9552 -3812 -8264 -2788
rect -8200 -3812 -8180 -2788
rect -9552 -3840 -8180 -3812
rect -7940 -2788 -6568 -2760
rect -7940 -3812 -6652 -2788
rect -6588 -3812 -6568 -2788
rect -7940 -3840 -6568 -3812
rect -6328 -2788 -4956 -2760
rect -6328 -3812 -5040 -2788
rect -4976 -3812 -4956 -2788
rect -6328 -3840 -4956 -3812
rect -4716 -2788 -3344 -2760
rect -4716 -3812 -3428 -2788
rect -3364 -3812 -3344 -2788
rect -4716 -3840 -3344 -3812
rect -3104 -2788 -1732 -2760
rect -3104 -3812 -1816 -2788
rect -1752 -3812 -1732 -2788
rect -3104 -3840 -1732 -3812
rect -1492 -2788 -120 -2760
rect -1492 -3812 -204 -2788
rect -140 -3812 -120 -2788
rect -1492 -3840 -120 -3812
rect 120 -2788 1492 -2760
rect 120 -3812 1408 -2788
rect 1472 -3812 1492 -2788
rect 120 -3840 1492 -3812
rect 1732 -2788 3104 -2760
rect 1732 -3812 3020 -2788
rect 3084 -3812 3104 -2788
rect 1732 -3840 3104 -3812
rect 3344 -2788 4716 -2760
rect 3344 -3812 4632 -2788
rect 4696 -3812 4716 -2788
rect 3344 -3840 4716 -3812
rect 4956 -2788 6328 -2760
rect 4956 -3812 6244 -2788
rect 6308 -3812 6328 -2788
rect 4956 -3840 6328 -3812
rect 6568 -2788 7940 -2760
rect 6568 -3812 7856 -2788
rect 7920 -3812 7940 -2788
rect 6568 -3840 7940 -3812
rect 8180 -2788 9552 -2760
rect 8180 -3812 9468 -2788
rect 9532 -3812 9552 -2788
rect 8180 -3840 9552 -3812
rect 9792 -2788 11164 -2760
rect 9792 -3812 11080 -2788
rect 11144 -3812 11164 -2788
rect 9792 -3840 11164 -3812
rect 11404 -2788 12776 -2760
rect 11404 -3812 12692 -2788
rect 12756 -3812 12776 -2788
rect 11404 -3840 12776 -3812
rect -12776 -4108 -11404 -4080
rect -12776 -5132 -11488 -4108
rect -11424 -5132 -11404 -4108
rect -12776 -5160 -11404 -5132
rect -11164 -4108 -9792 -4080
rect -11164 -5132 -9876 -4108
rect -9812 -5132 -9792 -4108
rect -11164 -5160 -9792 -5132
rect -9552 -4108 -8180 -4080
rect -9552 -5132 -8264 -4108
rect -8200 -5132 -8180 -4108
rect -9552 -5160 -8180 -5132
rect -7940 -4108 -6568 -4080
rect -7940 -5132 -6652 -4108
rect -6588 -5132 -6568 -4108
rect -7940 -5160 -6568 -5132
rect -6328 -4108 -4956 -4080
rect -6328 -5132 -5040 -4108
rect -4976 -5132 -4956 -4108
rect -6328 -5160 -4956 -5132
rect -4716 -4108 -3344 -4080
rect -4716 -5132 -3428 -4108
rect -3364 -5132 -3344 -4108
rect -4716 -5160 -3344 -5132
rect -3104 -4108 -1732 -4080
rect -3104 -5132 -1816 -4108
rect -1752 -5132 -1732 -4108
rect -3104 -5160 -1732 -5132
rect -1492 -4108 -120 -4080
rect -1492 -5132 -204 -4108
rect -140 -5132 -120 -4108
rect -1492 -5160 -120 -5132
rect 120 -4108 1492 -4080
rect 120 -5132 1408 -4108
rect 1472 -5132 1492 -4108
rect 120 -5160 1492 -5132
rect 1732 -4108 3104 -4080
rect 1732 -5132 3020 -4108
rect 3084 -5132 3104 -4108
rect 1732 -5160 3104 -5132
rect 3344 -4108 4716 -4080
rect 3344 -5132 4632 -4108
rect 4696 -5132 4716 -4108
rect 3344 -5160 4716 -5132
rect 4956 -4108 6328 -4080
rect 4956 -5132 6244 -4108
rect 6308 -5132 6328 -4108
rect 4956 -5160 6328 -5132
rect 6568 -4108 7940 -4080
rect 6568 -5132 7856 -4108
rect 7920 -5132 7940 -4108
rect 6568 -5160 7940 -5132
rect 8180 -4108 9552 -4080
rect 8180 -5132 9468 -4108
rect 9532 -5132 9552 -4108
rect 8180 -5160 9552 -5132
rect 9792 -4108 11164 -4080
rect 9792 -5132 11080 -4108
rect 11144 -5132 11164 -4108
rect 9792 -5160 11164 -5132
rect 11404 -4108 12776 -4080
rect 11404 -5132 12692 -4108
rect 12756 -5132 12776 -4108
rect 11404 -5160 12776 -5132
<< via3 >>
rect -11488 4108 -11424 5132
rect -9876 4108 -9812 5132
rect -8264 4108 -8200 5132
rect -6652 4108 -6588 5132
rect -5040 4108 -4976 5132
rect -3428 4108 -3364 5132
rect -1816 4108 -1752 5132
rect -204 4108 -140 5132
rect 1408 4108 1472 5132
rect 3020 4108 3084 5132
rect 4632 4108 4696 5132
rect 6244 4108 6308 5132
rect 7856 4108 7920 5132
rect 9468 4108 9532 5132
rect 11080 4108 11144 5132
rect 12692 4108 12756 5132
rect -11488 2788 -11424 3812
rect -9876 2788 -9812 3812
rect -8264 2788 -8200 3812
rect -6652 2788 -6588 3812
rect -5040 2788 -4976 3812
rect -3428 2788 -3364 3812
rect -1816 2788 -1752 3812
rect -204 2788 -140 3812
rect 1408 2788 1472 3812
rect 3020 2788 3084 3812
rect 4632 2788 4696 3812
rect 6244 2788 6308 3812
rect 7856 2788 7920 3812
rect 9468 2788 9532 3812
rect 11080 2788 11144 3812
rect 12692 2788 12756 3812
rect -11488 1468 -11424 2492
rect -9876 1468 -9812 2492
rect -8264 1468 -8200 2492
rect -6652 1468 -6588 2492
rect -5040 1468 -4976 2492
rect -3428 1468 -3364 2492
rect -1816 1468 -1752 2492
rect -204 1468 -140 2492
rect 1408 1468 1472 2492
rect 3020 1468 3084 2492
rect 4632 1468 4696 2492
rect 6244 1468 6308 2492
rect 7856 1468 7920 2492
rect 9468 1468 9532 2492
rect 11080 1468 11144 2492
rect 12692 1468 12756 2492
rect -11488 148 -11424 1172
rect -9876 148 -9812 1172
rect -8264 148 -8200 1172
rect -6652 148 -6588 1172
rect -5040 148 -4976 1172
rect -3428 148 -3364 1172
rect -1816 148 -1752 1172
rect -204 148 -140 1172
rect 1408 148 1472 1172
rect 3020 148 3084 1172
rect 4632 148 4696 1172
rect 6244 148 6308 1172
rect 7856 148 7920 1172
rect 9468 148 9532 1172
rect 11080 148 11144 1172
rect 12692 148 12756 1172
rect -11488 -1172 -11424 -148
rect -9876 -1172 -9812 -148
rect -8264 -1172 -8200 -148
rect -6652 -1172 -6588 -148
rect -5040 -1172 -4976 -148
rect -3428 -1172 -3364 -148
rect -1816 -1172 -1752 -148
rect -204 -1172 -140 -148
rect 1408 -1172 1472 -148
rect 3020 -1172 3084 -148
rect 4632 -1172 4696 -148
rect 6244 -1172 6308 -148
rect 7856 -1172 7920 -148
rect 9468 -1172 9532 -148
rect 11080 -1172 11144 -148
rect 12692 -1172 12756 -148
rect -11488 -2492 -11424 -1468
rect -9876 -2492 -9812 -1468
rect -8264 -2492 -8200 -1468
rect -6652 -2492 -6588 -1468
rect -5040 -2492 -4976 -1468
rect -3428 -2492 -3364 -1468
rect -1816 -2492 -1752 -1468
rect -204 -2492 -140 -1468
rect 1408 -2492 1472 -1468
rect 3020 -2492 3084 -1468
rect 4632 -2492 4696 -1468
rect 6244 -2492 6308 -1468
rect 7856 -2492 7920 -1468
rect 9468 -2492 9532 -1468
rect 11080 -2492 11144 -1468
rect 12692 -2492 12756 -1468
rect -11488 -3812 -11424 -2788
rect -9876 -3812 -9812 -2788
rect -8264 -3812 -8200 -2788
rect -6652 -3812 -6588 -2788
rect -5040 -3812 -4976 -2788
rect -3428 -3812 -3364 -2788
rect -1816 -3812 -1752 -2788
rect -204 -3812 -140 -2788
rect 1408 -3812 1472 -2788
rect 3020 -3812 3084 -2788
rect 4632 -3812 4696 -2788
rect 6244 -3812 6308 -2788
rect 7856 -3812 7920 -2788
rect 9468 -3812 9532 -2788
rect 11080 -3812 11144 -2788
rect 12692 -3812 12756 -2788
rect -11488 -5132 -11424 -4108
rect -9876 -5132 -9812 -4108
rect -8264 -5132 -8200 -4108
rect -6652 -5132 -6588 -4108
rect -5040 -5132 -4976 -4108
rect -3428 -5132 -3364 -4108
rect -1816 -5132 -1752 -4108
rect -204 -5132 -140 -4108
rect 1408 -5132 1472 -4108
rect 3020 -5132 3084 -4108
rect 4632 -5132 4696 -4108
rect 6244 -5132 6308 -4108
rect 7856 -5132 7920 -4108
rect 9468 -5132 9532 -4108
rect 11080 -5132 11144 -4108
rect 12692 -5132 12756 -4108
<< mimcap >>
rect -12736 5080 -11736 5120
rect -12736 4160 -12696 5080
rect -11776 4160 -11736 5080
rect -12736 4120 -11736 4160
rect -11124 5080 -10124 5120
rect -11124 4160 -11084 5080
rect -10164 4160 -10124 5080
rect -11124 4120 -10124 4160
rect -9512 5080 -8512 5120
rect -9512 4160 -9472 5080
rect -8552 4160 -8512 5080
rect -9512 4120 -8512 4160
rect -7900 5080 -6900 5120
rect -7900 4160 -7860 5080
rect -6940 4160 -6900 5080
rect -7900 4120 -6900 4160
rect -6288 5080 -5288 5120
rect -6288 4160 -6248 5080
rect -5328 4160 -5288 5080
rect -6288 4120 -5288 4160
rect -4676 5080 -3676 5120
rect -4676 4160 -4636 5080
rect -3716 4160 -3676 5080
rect -4676 4120 -3676 4160
rect -3064 5080 -2064 5120
rect -3064 4160 -3024 5080
rect -2104 4160 -2064 5080
rect -3064 4120 -2064 4160
rect -1452 5080 -452 5120
rect -1452 4160 -1412 5080
rect -492 4160 -452 5080
rect -1452 4120 -452 4160
rect 160 5080 1160 5120
rect 160 4160 200 5080
rect 1120 4160 1160 5080
rect 160 4120 1160 4160
rect 1772 5080 2772 5120
rect 1772 4160 1812 5080
rect 2732 4160 2772 5080
rect 1772 4120 2772 4160
rect 3384 5080 4384 5120
rect 3384 4160 3424 5080
rect 4344 4160 4384 5080
rect 3384 4120 4384 4160
rect 4996 5080 5996 5120
rect 4996 4160 5036 5080
rect 5956 4160 5996 5080
rect 4996 4120 5996 4160
rect 6608 5080 7608 5120
rect 6608 4160 6648 5080
rect 7568 4160 7608 5080
rect 6608 4120 7608 4160
rect 8220 5080 9220 5120
rect 8220 4160 8260 5080
rect 9180 4160 9220 5080
rect 8220 4120 9220 4160
rect 9832 5080 10832 5120
rect 9832 4160 9872 5080
rect 10792 4160 10832 5080
rect 9832 4120 10832 4160
rect 11444 5080 12444 5120
rect 11444 4160 11484 5080
rect 12404 4160 12444 5080
rect 11444 4120 12444 4160
rect -12736 3760 -11736 3800
rect -12736 2840 -12696 3760
rect -11776 2840 -11736 3760
rect -12736 2800 -11736 2840
rect -11124 3760 -10124 3800
rect -11124 2840 -11084 3760
rect -10164 2840 -10124 3760
rect -11124 2800 -10124 2840
rect -9512 3760 -8512 3800
rect -9512 2840 -9472 3760
rect -8552 2840 -8512 3760
rect -9512 2800 -8512 2840
rect -7900 3760 -6900 3800
rect -7900 2840 -7860 3760
rect -6940 2840 -6900 3760
rect -7900 2800 -6900 2840
rect -6288 3760 -5288 3800
rect -6288 2840 -6248 3760
rect -5328 2840 -5288 3760
rect -6288 2800 -5288 2840
rect -4676 3760 -3676 3800
rect -4676 2840 -4636 3760
rect -3716 2840 -3676 3760
rect -4676 2800 -3676 2840
rect -3064 3760 -2064 3800
rect -3064 2840 -3024 3760
rect -2104 2840 -2064 3760
rect -3064 2800 -2064 2840
rect -1452 3760 -452 3800
rect -1452 2840 -1412 3760
rect -492 2840 -452 3760
rect -1452 2800 -452 2840
rect 160 3760 1160 3800
rect 160 2840 200 3760
rect 1120 2840 1160 3760
rect 160 2800 1160 2840
rect 1772 3760 2772 3800
rect 1772 2840 1812 3760
rect 2732 2840 2772 3760
rect 1772 2800 2772 2840
rect 3384 3760 4384 3800
rect 3384 2840 3424 3760
rect 4344 2840 4384 3760
rect 3384 2800 4384 2840
rect 4996 3760 5996 3800
rect 4996 2840 5036 3760
rect 5956 2840 5996 3760
rect 4996 2800 5996 2840
rect 6608 3760 7608 3800
rect 6608 2840 6648 3760
rect 7568 2840 7608 3760
rect 6608 2800 7608 2840
rect 8220 3760 9220 3800
rect 8220 2840 8260 3760
rect 9180 2840 9220 3760
rect 8220 2800 9220 2840
rect 9832 3760 10832 3800
rect 9832 2840 9872 3760
rect 10792 2840 10832 3760
rect 9832 2800 10832 2840
rect 11444 3760 12444 3800
rect 11444 2840 11484 3760
rect 12404 2840 12444 3760
rect 11444 2800 12444 2840
rect -12736 2440 -11736 2480
rect -12736 1520 -12696 2440
rect -11776 1520 -11736 2440
rect -12736 1480 -11736 1520
rect -11124 2440 -10124 2480
rect -11124 1520 -11084 2440
rect -10164 1520 -10124 2440
rect -11124 1480 -10124 1520
rect -9512 2440 -8512 2480
rect -9512 1520 -9472 2440
rect -8552 1520 -8512 2440
rect -9512 1480 -8512 1520
rect -7900 2440 -6900 2480
rect -7900 1520 -7860 2440
rect -6940 1520 -6900 2440
rect -7900 1480 -6900 1520
rect -6288 2440 -5288 2480
rect -6288 1520 -6248 2440
rect -5328 1520 -5288 2440
rect -6288 1480 -5288 1520
rect -4676 2440 -3676 2480
rect -4676 1520 -4636 2440
rect -3716 1520 -3676 2440
rect -4676 1480 -3676 1520
rect -3064 2440 -2064 2480
rect -3064 1520 -3024 2440
rect -2104 1520 -2064 2440
rect -3064 1480 -2064 1520
rect -1452 2440 -452 2480
rect -1452 1520 -1412 2440
rect -492 1520 -452 2440
rect -1452 1480 -452 1520
rect 160 2440 1160 2480
rect 160 1520 200 2440
rect 1120 1520 1160 2440
rect 160 1480 1160 1520
rect 1772 2440 2772 2480
rect 1772 1520 1812 2440
rect 2732 1520 2772 2440
rect 1772 1480 2772 1520
rect 3384 2440 4384 2480
rect 3384 1520 3424 2440
rect 4344 1520 4384 2440
rect 3384 1480 4384 1520
rect 4996 2440 5996 2480
rect 4996 1520 5036 2440
rect 5956 1520 5996 2440
rect 4996 1480 5996 1520
rect 6608 2440 7608 2480
rect 6608 1520 6648 2440
rect 7568 1520 7608 2440
rect 6608 1480 7608 1520
rect 8220 2440 9220 2480
rect 8220 1520 8260 2440
rect 9180 1520 9220 2440
rect 8220 1480 9220 1520
rect 9832 2440 10832 2480
rect 9832 1520 9872 2440
rect 10792 1520 10832 2440
rect 9832 1480 10832 1520
rect 11444 2440 12444 2480
rect 11444 1520 11484 2440
rect 12404 1520 12444 2440
rect 11444 1480 12444 1520
rect -12736 1120 -11736 1160
rect -12736 200 -12696 1120
rect -11776 200 -11736 1120
rect -12736 160 -11736 200
rect -11124 1120 -10124 1160
rect -11124 200 -11084 1120
rect -10164 200 -10124 1120
rect -11124 160 -10124 200
rect -9512 1120 -8512 1160
rect -9512 200 -9472 1120
rect -8552 200 -8512 1120
rect -9512 160 -8512 200
rect -7900 1120 -6900 1160
rect -7900 200 -7860 1120
rect -6940 200 -6900 1120
rect -7900 160 -6900 200
rect -6288 1120 -5288 1160
rect -6288 200 -6248 1120
rect -5328 200 -5288 1120
rect -6288 160 -5288 200
rect -4676 1120 -3676 1160
rect -4676 200 -4636 1120
rect -3716 200 -3676 1120
rect -4676 160 -3676 200
rect -3064 1120 -2064 1160
rect -3064 200 -3024 1120
rect -2104 200 -2064 1120
rect -3064 160 -2064 200
rect -1452 1120 -452 1160
rect -1452 200 -1412 1120
rect -492 200 -452 1120
rect -1452 160 -452 200
rect 160 1120 1160 1160
rect 160 200 200 1120
rect 1120 200 1160 1120
rect 160 160 1160 200
rect 1772 1120 2772 1160
rect 1772 200 1812 1120
rect 2732 200 2772 1120
rect 1772 160 2772 200
rect 3384 1120 4384 1160
rect 3384 200 3424 1120
rect 4344 200 4384 1120
rect 3384 160 4384 200
rect 4996 1120 5996 1160
rect 4996 200 5036 1120
rect 5956 200 5996 1120
rect 4996 160 5996 200
rect 6608 1120 7608 1160
rect 6608 200 6648 1120
rect 7568 200 7608 1120
rect 6608 160 7608 200
rect 8220 1120 9220 1160
rect 8220 200 8260 1120
rect 9180 200 9220 1120
rect 8220 160 9220 200
rect 9832 1120 10832 1160
rect 9832 200 9872 1120
rect 10792 200 10832 1120
rect 9832 160 10832 200
rect 11444 1120 12444 1160
rect 11444 200 11484 1120
rect 12404 200 12444 1120
rect 11444 160 12444 200
rect -12736 -200 -11736 -160
rect -12736 -1120 -12696 -200
rect -11776 -1120 -11736 -200
rect -12736 -1160 -11736 -1120
rect -11124 -200 -10124 -160
rect -11124 -1120 -11084 -200
rect -10164 -1120 -10124 -200
rect -11124 -1160 -10124 -1120
rect -9512 -200 -8512 -160
rect -9512 -1120 -9472 -200
rect -8552 -1120 -8512 -200
rect -9512 -1160 -8512 -1120
rect -7900 -200 -6900 -160
rect -7900 -1120 -7860 -200
rect -6940 -1120 -6900 -200
rect -7900 -1160 -6900 -1120
rect -6288 -200 -5288 -160
rect -6288 -1120 -6248 -200
rect -5328 -1120 -5288 -200
rect -6288 -1160 -5288 -1120
rect -4676 -200 -3676 -160
rect -4676 -1120 -4636 -200
rect -3716 -1120 -3676 -200
rect -4676 -1160 -3676 -1120
rect -3064 -200 -2064 -160
rect -3064 -1120 -3024 -200
rect -2104 -1120 -2064 -200
rect -3064 -1160 -2064 -1120
rect -1452 -200 -452 -160
rect -1452 -1120 -1412 -200
rect -492 -1120 -452 -200
rect -1452 -1160 -452 -1120
rect 160 -200 1160 -160
rect 160 -1120 200 -200
rect 1120 -1120 1160 -200
rect 160 -1160 1160 -1120
rect 1772 -200 2772 -160
rect 1772 -1120 1812 -200
rect 2732 -1120 2772 -200
rect 1772 -1160 2772 -1120
rect 3384 -200 4384 -160
rect 3384 -1120 3424 -200
rect 4344 -1120 4384 -200
rect 3384 -1160 4384 -1120
rect 4996 -200 5996 -160
rect 4996 -1120 5036 -200
rect 5956 -1120 5996 -200
rect 4996 -1160 5996 -1120
rect 6608 -200 7608 -160
rect 6608 -1120 6648 -200
rect 7568 -1120 7608 -200
rect 6608 -1160 7608 -1120
rect 8220 -200 9220 -160
rect 8220 -1120 8260 -200
rect 9180 -1120 9220 -200
rect 8220 -1160 9220 -1120
rect 9832 -200 10832 -160
rect 9832 -1120 9872 -200
rect 10792 -1120 10832 -200
rect 9832 -1160 10832 -1120
rect 11444 -200 12444 -160
rect 11444 -1120 11484 -200
rect 12404 -1120 12444 -200
rect 11444 -1160 12444 -1120
rect -12736 -1520 -11736 -1480
rect -12736 -2440 -12696 -1520
rect -11776 -2440 -11736 -1520
rect -12736 -2480 -11736 -2440
rect -11124 -1520 -10124 -1480
rect -11124 -2440 -11084 -1520
rect -10164 -2440 -10124 -1520
rect -11124 -2480 -10124 -2440
rect -9512 -1520 -8512 -1480
rect -9512 -2440 -9472 -1520
rect -8552 -2440 -8512 -1520
rect -9512 -2480 -8512 -2440
rect -7900 -1520 -6900 -1480
rect -7900 -2440 -7860 -1520
rect -6940 -2440 -6900 -1520
rect -7900 -2480 -6900 -2440
rect -6288 -1520 -5288 -1480
rect -6288 -2440 -6248 -1520
rect -5328 -2440 -5288 -1520
rect -6288 -2480 -5288 -2440
rect -4676 -1520 -3676 -1480
rect -4676 -2440 -4636 -1520
rect -3716 -2440 -3676 -1520
rect -4676 -2480 -3676 -2440
rect -3064 -1520 -2064 -1480
rect -3064 -2440 -3024 -1520
rect -2104 -2440 -2064 -1520
rect -3064 -2480 -2064 -2440
rect -1452 -1520 -452 -1480
rect -1452 -2440 -1412 -1520
rect -492 -2440 -452 -1520
rect -1452 -2480 -452 -2440
rect 160 -1520 1160 -1480
rect 160 -2440 200 -1520
rect 1120 -2440 1160 -1520
rect 160 -2480 1160 -2440
rect 1772 -1520 2772 -1480
rect 1772 -2440 1812 -1520
rect 2732 -2440 2772 -1520
rect 1772 -2480 2772 -2440
rect 3384 -1520 4384 -1480
rect 3384 -2440 3424 -1520
rect 4344 -2440 4384 -1520
rect 3384 -2480 4384 -2440
rect 4996 -1520 5996 -1480
rect 4996 -2440 5036 -1520
rect 5956 -2440 5996 -1520
rect 4996 -2480 5996 -2440
rect 6608 -1520 7608 -1480
rect 6608 -2440 6648 -1520
rect 7568 -2440 7608 -1520
rect 6608 -2480 7608 -2440
rect 8220 -1520 9220 -1480
rect 8220 -2440 8260 -1520
rect 9180 -2440 9220 -1520
rect 8220 -2480 9220 -2440
rect 9832 -1520 10832 -1480
rect 9832 -2440 9872 -1520
rect 10792 -2440 10832 -1520
rect 9832 -2480 10832 -2440
rect 11444 -1520 12444 -1480
rect 11444 -2440 11484 -1520
rect 12404 -2440 12444 -1520
rect 11444 -2480 12444 -2440
rect -12736 -2840 -11736 -2800
rect -12736 -3760 -12696 -2840
rect -11776 -3760 -11736 -2840
rect -12736 -3800 -11736 -3760
rect -11124 -2840 -10124 -2800
rect -11124 -3760 -11084 -2840
rect -10164 -3760 -10124 -2840
rect -11124 -3800 -10124 -3760
rect -9512 -2840 -8512 -2800
rect -9512 -3760 -9472 -2840
rect -8552 -3760 -8512 -2840
rect -9512 -3800 -8512 -3760
rect -7900 -2840 -6900 -2800
rect -7900 -3760 -7860 -2840
rect -6940 -3760 -6900 -2840
rect -7900 -3800 -6900 -3760
rect -6288 -2840 -5288 -2800
rect -6288 -3760 -6248 -2840
rect -5328 -3760 -5288 -2840
rect -6288 -3800 -5288 -3760
rect -4676 -2840 -3676 -2800
rect -4676 -3760 -4636 -2840
rect -3716 -3760 -3676 -2840
rect -4676 -3800 -3676 -3760
rect -3064 -2840 -2064 -2800
rect -3064 -3760 -3024 -2840
rect -2104 -3760 -2064 -2840
rect -3064 -3800 -2064 -3760
rect -1452 -2840 -452 -2800
rect -1452 -3760 -1412 -2840
rect -492 -3760 -452 -2840
rect -1452 -3800 -452 -3760
rect 160 -2840 1160 -2800
rect 160 -3760 200 -2840
rect 1120 -3760 1160 -2840
rect 160 -3800 1160 -3760
rect 1772 -2840 2772 -2800
rect 1772 -3760 1812 -2840
rect 2732 -3760 2772 -2840
rect 1772 -3800 2772 -3760
rect 3384 -2840 4384 -2800
rect 3384 -3760 3424 -2840
rect 4344 -3760 4384 -2840
rect 3384 -3800 4384 -3760
rect 4996 -2840 5996 -2800
rect 4996 -3760 5036 -2840
rect 5956 -3760 5996 -2840
rect 4996 -3800 5996 -3760
rect 6608 -2840 7608 -2800
rect 6608 -3760 6648 -2840
rect 7568 -3760 7608 -2840
rect 6608 -3800 7608 -3760
rect 8220 -2840 9220 -2800
rect 8220 -3760 8260 -2840
rect 9180 -3760 9220 -2840
rect 8220 -3800 9220 -3760
rect 9832 -2840 10832 -2800
rect 9832 -3760 9872 -2840
rect 10792 -3760 10832 -2840
rect 9832 -3800 10832 -3760
rect 11444 -2840 12444 -2800
rect 11444 -3760 11484 -2840
rect 12404 -3760 12444 -2840
rect 11444 -3800 12444 -3760
rect -12736 -4160 -11736 -4120
rect -12736 -5080 -12696 -4160
rect -11776 -5080 -11736 -4160
rect -12736 -5120 -11736 -5080
rect -11124 -4160 -10124 -4120
rect -11124 -5080 -11084 -4160
rect -10164 -5080 -10124 -4160
rect -11124 -5120 -10124 -5080
rect -9512 -4160 -8512 -4120
rect -9512 -5080 -9472 -4160
rect -8552 -5080 -8512 -4160
rect -9512 -5120 -8512 -5080
rect -7900 -4160 -6900 -4120
rect -7900 -5080 -7860 -4160
rect -6940 -5080 -6900 -4160
rect -7900 -5120 -6900 -5080
rect -6288 -4160 -5288 -4120
rect -6288 -5080 -6248 -4160
rect -5328 -5080 -5288 -4160
rect -6288 -5120 -5288 -5080
rect -4676 -4160 -3676 -4120
rect -4676 -5080 -4636 -4160
rect -3716 -5080 -3676 -4160
rect -4676 -5120 -3676 -5080
rect -3064 -4160 -2064 -4120
rect -3064 -5080 -3024 -4160
rect -2104 -5080 -2064 -4160
rect -3064 -5120 -2064 -5080
rect -1452 -4160 -452 -4120
rect -1452 -5080 -1412 -4160
rect -492 -5080 -452 -4160
rect -1452 -5120 -452 -5080
rect 160 -4160 1160 -4120
rect 160 -5080 200 -4160
rect 1120 -5080 1160 -4160
rect 160 -5120 1160 -5080
rect 1772 -4160 2772 -4120
rect 1772 -5080 1812 -4160
rect 2732 -5080 2772 -4160
rect 1772 -5120 2772 -5080
rect 3384 -4160 4384 -4120
rect 3384 -5080 3424 -4160
rect 4344 -5080 4384 -4160
rect 3384 -5120 4384 -5080
rect 4996 -4160 5996 -4120
rect 4996 -5080 5036 -4160
rect 5956 -5080 5996 -4160
rect 4996 -5120 5996 -5080
rect 6608 -4160 7608 -4120
rect 6608 -5080 6648 -4160
rect 7568 -5080 7608 -4160
rect 6608 -5120 7608 -5080
rect 8220 -4160 9220 -4120
rect 8220 -5080 8260 -4160
rect 9180 -5080 9220 -4160
rect 8220 -5120 9220 -5080
rect 9832 -4160 10832 -4120
rect 9832 -5080 9872 -4160
rect 10792 -5080 10832 -4160
rect 9832 -5120 10832 -5080
rect 11444 -4160 12444 -4120
rect 11444 -5080 11484 -4160
rect 12404 -5080 12444 -4160
rect 11444 -5120 12444 -5080
<< mimcapcontact >>
rect -12696 4160 -11776 5080
rect -11084 4160 -10164 5080
rect -9472 4160 -8552 5080
rect -7860 4160 -6940 5080
rect -6248 4160 -5328 5080
rect -4636 4160 -3716 5080
rect -3024 4160 -2104 5080
rect -1412 4160 -492 5080
rect 200 4160 1120 5080
rect 1812 4160 2732 5080
rect 3424 4160 4344 5080
rect 5036 4160 5956 5080
rect 6648 4160 7568 5080
rect 8260 4160 9180 5080
rect 9872 4160 10792 5080
rect 11484 4160 12404 5080
rect -12696 2840 -11776 3760
rect -11084 2840 -10164 3760
rect -9472 2840 -8552 3760
rect -7860 2840 -6940 3760
rect -6248 2840 -5328 3760
rect -4636 2840 -3716 3760
rect -3024 2840 -2104 3760
rect -1412 2840 -492 3760
rect 200 2840 1120 3760
rect 1812 2840 2732 3760
rect 3424 2840 4344 3760
rect 5036 2840 5956 3760
rect 6648 2840 7568 3760
rect 8260 2840 9180 3760
rect 9872 2840 10792 3760
rect 11484 2840 12404 3760
rect -12696 1520 -11776 2440
rect -11084 1520 -10164 2440
rect -9472 1520 -8552 2440
rect -7860 1520 -6940 2440
rect -6248 1520 -5328 2440
rect -4636 1520 -3716 2440
rect -3024 1520 -2104 2440
rect -1412 1520 -492 2440
rect 200 1520 1120 2440
rect 1812 1520 2732 2440
rect 3424 1520 4344 2440
rect 5036 1520 5956 2440
rect 6648 1520 7568 2440
rect 8260 1520 9180 2440
rect 9872 1520 10792 2440
rect 11484 1520 12404 2440
rect -12696 200 -11776 1120
rect -11084 200 -10164 1120
rect -9472 200 -8552 1120
rect -7860 200 -6940 1120
rect -6248 200 -5328 1120
rect -4636 200 -3716 1120
rect -3024 200 -2104 1120
rect -1412 200 -492 1120
rect 200 200 1120 1120
rect 1812 200 2732 1120
rect 3424 200 4344 1120
rect 5036 200 5956 1120
rect 6648 200 7568 1120
rect 8260 200 9180 1120
rect 9872 200 10792 1120
rect 11484 200 12404 1120
rect -12696 -1120 -11776 -200
rect -11084 -1120 -10164 -200
rect -9472 -1120 -8552 -200
rect -7860 -1120 -6940 -200
rect -6248 -1120 -5328 -200
rect -4636 -1120 -3716 -200
rect -3024 -1120 -2104 -200
rect -1412 -1120 -492 -200
rect 200 -1120 1120 -200
rect 1812 -1120 2732 -200
rect 3424 -1120 4344 -200
rect 5036 -1120 5956 -200
rect 6648 -1120 7568 -200
rect 8260 -1120 9180 -200
rect 9872 -1120 10792 -200
rect 11484 -1120 12404 -200
rect -12696 -2440 -11776 -1520
rect -11084 -2440 -10164 -1520
rect -9472 -2440 -8552 -1520
rect -7860 -2440 -6940 -1520
rect -6248 -2440 -5328 -1520
rect -4636 -2440 -3716 -1520
rect -3024 -2440 -2104 -1520
rect -1412 -2440 -492 -1520
rect 200 -2440 1120 -1520
rect 1812 -2440 2732 -1520
rect 3424 -2440 4344 -1520
rect 5036 -2440 5956 -1520
rect 6648 -2440 7568 -1520
rect 8260 -2440 9180 -1520
rect 9872 -2440 10792 -1520
rect 11484 -2440 12404 -1520
rect -12696 -3760 -11776 -2840
rect -11084 -3760 -10164 -2840
rect -9472 -3760 -8552 -2840
rect -7860 -3760 -6940 -2840
rect -6248 -3760 -5328 -2840
rect -4636 -3760 -3716 -2840
rect -3024 -3760 -2104 -2840
rect -1412 -3760 -492 -2840
rect 200 -3760 1120 -2840
rect 1812 -3760 2732 -2840
rect 3424 -3760 4344 -2840
rect 5036 -3760 5956 -2840
rect 6648 -3760 7568 -2840
rect 8260 -3760 9180 -2840
rect 9872 -3760 10792 -2840
rect 11484 -3760 12404 -2840
rect -12696 -5080 -11776 -4160
rect -11084 -5080 -10164 -4160
rect -9472 -5080 -8552 -4160
rect -7860 -5080 -6940 -4160
rect -6248 -5080 -5328 -4160
rect -4636 -5080 -3716 -4160
rect -3024 -5080 -2104 -4160
rect -1412 -5080 -492 -4160
rect 200 -5080 1120 -4160
rect 1812 -5080 2732 -4160
rect 3424 -5080 4344 -4160
rect 5036 -5080 5956 -4160
rect 6648 -5080 7568 -4160
rect 8260 -5080 9180 -4160
rect 9872 -5080 10792 -4160
rect 11484 -5080 12404 -4160
<< metal4 >>
rect -12288 5081 -12184 5280
rect -11508 5132 -11404 5280
rect -12697 5080 -11775 5081
rect -12697 4160 -12696 5080
rect -11776 4160 -11775 5080
rect -12697 4159 -11775 4160
rect -12288 3761 -12184 4159
rect -11508 4108 -11488 5132
rect -11424 4108 -11404 5132
rect -10676 5081 -10572 5280
rect -9896 5132 -9792 5280
rect -11085 5080 -10163 5081
rect -11085 4160 -11084 5080
rect -10164 4160 -10163 5080
rect -11085 4159 -10163 4160
rect -11508 3812 -11404 4108
rect -12697 3760 -11775 3761
rect -12697 2840 -12696 3760
rect -11776 2840 -11775 3760
rect -12697 2839 -11775 2840
rect -12288 2441 -12184 2839
rect -11508 2788 -11488 3812
rect -11424 2788 -11404 3812
rect -10676 3761 -10572 4159
rect -9896 4108 -9876 5132
rect -9812 4108 -9792 5132
rect -9064 5081 -8960 5280
rect -8284 5132 -8180 5280
rect -9473 5080 -8551 5081
rect -9473 4160 -9472 5080
rect -8552 4160 -8551 5080
rect -9473 4159 -8551 4160
rect -9896 3812 -9792 4108
rect -11085 3760 -10163 3761
rect -11085 2840 -11084 3760
rect -10164 2840 -10163 3760
rect -11085 2839 -10163 2840
rect -11508 2492 -11404 2788
rect -12697 2440 -11775 2441
rect -12697 1520 -12696 2440
rect -11776 1520 -11775 2440
rect -12697 1519 -11775 1520
rect -12288 1121 -12184 1519
rect -11508 1468 -11488 2492
rect -11424 1468 -11404 2492
rect -10676 2441 -10572 2839
rect -9896 2788 -9876 3812
rect -9812 2788 -9792 3812
rect -9064 3761 -8960 4159
rect -8284 4108 -8264 5132
rect -8200 4108 -8180 5132
rect -7452 5081 -7348 5280
rect -6672 5132 -6568 5280
rect -7861 5080 -6939 5081
rect -7861 4160 -7860 5080
rect -6940 4160 -6939 5080
rect -7861 4159 -6939 4160
rect -8284 3812 -8180 4108
rect -9473 3760 -8551 3761
rect -9473 2840 -9472 3760
rect -8552 2840 -8551 3760
rect -9473 2839 -8551 2840
rect -9896 2492 -9792 2788
rect -11085 2440 -10163 2441
rect -11085 1520 -11084 2440
rect -10164 1520 -10163 2440
rect -11085 1519 -10163 1520
rect -11508 1172 -11404 1468
rect -12697 1120 -11775 1121
rect -12697 200 -12696 1120
rect -11776 200 -11775 1120
rect -12697 199 -11775 200
rect -12288 -199 -12184 199
rect -11508 148 -11488 1172
rect -11424 148 -11404 1172
rect -10676 1121 -10572 1519
rect -9896 1468 -9876 2492
rect -9812 1468 -9792 2492
rect -9064 2441 -8960 2839
rect -8284 2788 -8264 3812
rect -8200 2788 -8180 3812
rect -7452 3761 -7348 4159
rect -6672 4108 -6652 5132
rect -6588 4108 -6568 5132
rect -5840 5081 -5736 5280
rect -5060 5132 -4956 5280
rect -6249 5080 -5327 5081
rect -6249 4160 -6248 5080
rect -5328 4160 -5327 5080
rect -6249 4159 -5327 4160
rect -6672 3812 -6568 4108
rect -7861 3760 -6939 3761
rect -7861 2840 -7860 3760
rect -6940 2840 -6939 3760
rect -7861 2839 -6939 2840
rect -8284 2492 -8180 2788
rect -9473 2440 -8551 2441
rect -9473 1520 -9472 2440
rect -8552 1520 -8551 2440
rect -9473 1519 -8551 1520
rect -9896 1172 -9792 1468
rect -11085 1120 -10163 1121
rect -11085 200 -11084 1120
rect -10164 200 -10163 1120
rect -11085 199 -10163 200
rect -11508 -148 -11404 148
rect -12697 -200 -11775 -199
rect -12697 -1120 -12696 -200
rect -11776 -1120 -11775 -200
rect -12697 -1121 -11775 -1120
rect -12288 -1519 -12184 -1121
rect -11508 -1172 -11488 -148
rect -11424 -1172 -11404 -148
rect -10676 -199 -10572 199
rect -9896 148 -9876 1172
rect -9812 148 -9792 1172
rect -9064 1121 -8960 1519
rect -8284 1468 -8264 2492
rect -8200 1468 -8180 2492
rect -7452 2441 -7348 2839
rect -6672 2788 -6652 3812
rect -6588 2788 -6568 3812
rect -5840 3761 -5736 4159
rect -5060 4108 -5040 5132
rect -4976 4108 -4956 5132
rect -4228 5081 -4124 5280
rect -3448 5132 -3344 5280
rect -4637 5080 -3715 5081
rect -4637 4160 -4636 5080
rect -3716 4160 -3715 5080
rect -4637 4159 -3715 4160
rect -5060 3812 -4956 4108
rect -6249 3760 -5327 3761
rect -6249 2840 -6248 3760
rect -5328 2840 -5327 3760
rect -6249 2839 -5327 2840
rect -6672 2492 -6568 2788
rect -7861 2440 -6939 2441
rect -7861 1520 -7860 2440
rect -6940 1520 -6939 2440
rect -7861 1519 -6939 1520
rect -8284 1172 -8180 1468
rect -9473 1120 -8551 1121
rect -9473 200 -9472 1120
rect -8552 200 -8551 1120
rect -9473 199 -8551 200
rect -9896 -148 -9792 148
rect -11085 -200 -10163 -199
rect -11085 -1120 -11084 -200
rect -10164 -1120 -10163 -200
rect -11085 -1121 -10163 -1120
rect -11508 -1468 -11404 -1172
rect -12697 -1520 -11775 -1519
rect -12697 -2440 -12696 -1520
rect -11776 -2440 -11775 -1520
rect -12697 -2441 -11775 -2440
rect -12288 -2839 -12184 -2441
rect -11508 -2492 -11488 -1468
rect -11424 -2492 -11404 -1468
rect -10676 -1519 -10572 -1121
rect -9896 -1172 -9876 -148
rect -9812 -1172 -9792 -148
rect -9064 -199 -8960 199
rect -8284 148 -8264 1172
rect -8200 148 -8180 1172
rect -7452 1121 -7348 1519
rect -6672 1468 -6652 2492
rect -6588 1468 -6568 2492
rect -5840 2441 -5736 2839
rect -5060 2788 -5040 3812
rect -4976 2788 -4956 3812
rect -4228 3761 -4124 4159
rect -3448 4108 -3428 5132
rect -3364 4108 -3344 5132
rect -2616 5081 -2512 5280
rect -1836 5132 -1732 5280
rect -3025 5080 -2103 5081
rect -3025 4160 -3024 5080
rect -2104 4160 -2103 5080
rect -3025 4159 -2103 4160
rect -3448 3812 -3344 4108
rect -4637 3760 -3715 3761
rect -4637 2840 -4636 3760
rect -3716 2840 -3715 3760
rect -4637 2839 -3715 2840
rect -5060 2492 -4956 2788
rect -6249 2440 -5327 2441
rect -6249 1520 -6248 2440
rect -5328 1520 -5327 2440
rect -6249 1519 -5327 1520
rect -6672 1172 -6568 1468
rect -7861 1120 -6939 1121
rect -7861 200 -7860 1120
rect -6940 200 -6939 1120
rect -7861 199 -6939 200
rect -8284 -148 -8180 148
rect -9473 -200 -8551 -199
rect -9473 -1120 -9472 -200
rect -8552 -1120 -8551 -200
rect -9473 -1121 -8551 -1120
rect -9896 -1468 -9792 -1172
rect -11085 -1520 -10163 -1519
rect -11085 -2440 -11084 -1520
rect -10164 -2440 -10163 -1520
rect -11085 -2441 -10163 -2440
rect -11508 -2788 -11404 -2492
rect -12697 -2840 -11775 -2839
rect -12697 -3760 -12696 -2840
rect -11776 -3760 -11775 -2840
rect -12697 -3761 -11775 -3760
rect -12288 -4159 -12184 -3761
rect -11508 -3812 -11488 -2788
rect -11424 -3812 -11404 -2788
rect -10676 -2839 -10572 -2441
rect -9896 -2492 -9876 -1468
rect -9812 -2492 -9792 -1468
rect -9064 -1519 -8960 -1121
rect -8284 -1172 -8264 -148
rect -8200 -1172 -8180 -148
rect -7452 -199 -7348 199
rect -6672 148 -6652 1172
rect -6588 148 -6568 1172
rect -5840 1121 -5736 1519
rect -5060 1468 -5040 2492
rect -4976 1468 -4956 2492
rect -4228 2441 -4124 2839
rect -3448 2788 -3428 3812
rect -3364 2788 -3344 3812
rect -2616 3761 -2512 4159
rect -1836 4108 -1816 5132
rect -1752 4108 -1732 5132
rect -1004 5081 -900 5280
rect -224 5132 -120 5280
rect -1413 5080 -491 5081
rect -1413 4160 -1412 5080
rect -492 4160 -491 5080
rect -1413 4159 -491 4160
rect -1836 3812 -1732 4108
rect -3025 3760 -2103 3761
rect -3025 2840 -3024 3760
rect -2104 2840 -2103 3760
rect -3025 2839 -2103 2840
rect -3448 2492 -3344 2788
rect -4637 2440 -3715 2441
rect -4637 1520 -4636 2440
rect -3716 1520 -3715 2440
rect -4637 1519 -3715 1520
rect -5060 1172 -4956 1468
rect -6249 1120 -5327 1121
rect -6249 200 -6248 1120
rect -5328 200 -5327 1120
rect -6249 199 -5327 200
rect -6672 -148 -6568 148
rect -7861 -200 -6939 -199
rect -7861 -1120 -7860 -200
rect -6940 -1120 -6939 -200
rect -7861 -1121 -6939 -1120
rect -8284 -1468 -8180 -1172
rect -9473 -1520 -8551 -1519
rect -9473 -2440 -9472 -1520
rect -8552 -2440 -8551 -1520
rect -9473 -2441 -8551 -2440
rect -9896 -2788 -9792 -2492
rect -11085 -2840 -10163 -2839
rect -11085 -3760 -11084 -2840
rect -10164 -3760 -10163 -2840
rect -11085 -3761 -10163 -3760
rect -11508 -4108 -11404 -3812
rect -12697 -4160 -11775 -4159
rect -12697 -5080 -12696 -4160
rect -11776 -5080 -11775 -4160
rect -12697 -5081 -11775 -5080
rect -12288 -5280 -12184 -5081
rect -11508 -5132 -11488 -4108
rect -11424 -5132 -11404 -4108
rect -10676 -4159 -10572 -3761
rect -9896 -3812 -9876 -2788
rect -9812 -3812 -9792 -2788
rect -9064 -2839 -8960 -2441
rect -8284 -2492 -8264 -1468
rect -8200 -2492 -8180 -1468
rect -7452 -1519 -7348 -1121
rect -6672 -1172 -6652 -148
rect -6588 -1172 -6568 -148
rect -5840 -199 -5736 199
rect -5060 148 -5040 1172
rect -4976 148 -4956 1172
rect -4228 1121 -4124 1519
rect -3448 1468 -3428 2492
rect -3364 1468 -3344 2492
rect -2616 2441 -2512 2839
rect -1836 2788 -1816 3812
rect -1752 2788 -1732 3812
rect -1004 3761 -900 4159
rect -224 4108 -204 5132
rect -140 4108 -120 5132
rect 608 5081 712 5280
rect 1388 5132 1492 5280
rect 199 5080 1121 5081
rect 199 4160 200 5080
rect 1120 4160 1121 5080
rect 199 4159 1121 4160
rect -224 3812 -120 4108
rect -1413 3760 -491 3761
rect -1413 2840 -1412 3760
rect -492 2840 -491 3760
rect -1413 2839 -491 2840
rect -1836 2492 -1732 2788
rect -3025 2440 -2103 2441
rect -3025 1520 -3024 2440
rect -2104 1520 -2103 2440
rect -3025 1519 -2103 1520
rect -3448 1172 -3344 1468
rect -4637 1120 -3715 1121
rect -4637 200 -4636 1120
rect -3716 200 -3715 1120
rect -4637 199 -3715 200
rect -5060 -148 -4956 148
rect -6249 -200 -5327 -199
rect -6249 -1120 -6248 -200
rect -5328 -1120 -5327 -200
rect -6249 -1121 -5327 -1120
rect -6672 -1468 -6568 -1172
rect -7861 -1520 -6939 -1519
rect -7861 -2440 -7860 -1520
rect -6940 -2440 -6939 -1520
rect -7861 -2441 -6939 -2440
rect -8284 -2788 -8180 -2492
rect -9473 -2840 -8551 -2839
rect -9473 -3760 -9472 -2840
rect -8552 -3760 -8551 -2840
rect -9473 -3761 -8551 -3760
rect -9896 -4108 -9792 -3812
rect -11085 -4160 -10163 -4159
rect -11085 -5080 -11084 -4160
rect -10164 -5080 -10163 -4160
rect -11085 -5081 -10163 -5080
rect -11508 -5280 -11404 -5132
rect -10676 -5280 -10572 -5081
rect -9896 -5132 -9876 -4108
rect -9812 -5132 -9792 -4108
rect -9064 -4159 -8960 -3761
rect -8284 -3812 -8264 -2788
rect -8200 -3812 -8180 -2788
rect -7452 -2839 -7348 -2441
rect -6672 -2492 -6652 -1468
rect -6588 -2492 -6568 -1468
rect -5840 -1519 -5736 -1121
rect -5060 -1172 -5040 -148
rect -4976 -1172 -4956 -148
rect -4228 -199 -4124 199
rect -3448 148 -3428 1172
rect -3364 148 -3344 1172
rect -2616 1121 -2512 1519
rect -1836 1468 -1816 2492
rect -1752 1468 -1732 2492
rect -1004 2441 -900 2839
rect -224 2788 -204 3812
rect -140 2788 -120 3812
rect 608 3761 712 4159
rect 1388 4108 1408 5132
rect 1472 4108 1492 5132
rect 2220 5081 2324 5280
rect 3000 5132 3104 5280
rect 1811 5080 2733 5081
rect 1811 4160 1812 5080
rect 2732 4160 2733 5080
rect 1811 4159 2733 4160
rect 1388 3812 1492 4108
rect 199 3760 1121 3761
rect 199 2840 200 3760
rect 1120 2840 1121 3760
rect 199 2839 1121 2840
rect -224 2492 -120 2788
rect -1413 2440 -491 2441
rect -1413 1520 -1412 2440
rect -492 1520 -491 2440
rect -1413 1519 -491 1520
rect -1836 1172 -1732 1468
rect -3025 1120 -2103 1121
rect -3025 200 -3024 1120
rect -2104 200 -2103 1120
rect -3025 199 -2103 200
rect -3448 -148 -3344 148
rect -4637 -200 -3715 -199
rect -4637 -1120 -4636 -200
rect -3716 -1120 -3715 -200
rect -4637 -1121 -3715 -1120
rect -5060 -1468 -4956 -1172
rect -6249 -1520 -5327 -1519
rect -6249 -2440 -6248 -1520
rect -5328 -2440 -5327 -1520
rect -6249 -2441 -5327 -2440
rect -6672 -2788 -6568 -2492
rect -7861 -2840 -6939 -2839
rect -7861 -3760 -7860 -2840
rect -6940 -3760 -6939 -2840
rect -7861 -3761 -6939 -3760
rect -8284 -4108 -8180 -3812
rect -9473 -4160 -8551 -4159
rect -9473 -5080 -9472 -4160
rect -8552 -5080 -8551 -4160
rect -9473 -5081 -8551 -5080
rect -9896 -5280 -9792 -5132
rect -9064 -5280 -8960 -5081
rect -8284 -5132 -8264 -4108
rect -8200 -5132 -8180 -4108
rect -7452 -4159 -7348 -3761
rect -6672 -3812 -6652 -2788
rect -6588 -3812 -6568 -2788
rect -5840 -2839 -5736 -2441
rect -5060 -2492 -5040 -1468
rect -4976 -2492 -4956 -1468
rect -4228 -1519 -4124 -1121
rect -3448 -1172 -3428 -148
rect -3364 -1172 -3344 -148
rect -2616 -199 -2512 199
rect -1836 148 -1816 1172
rect -1752 148 -1732 1172
rect -1004 1121 -900 1519
rect -224 1468 -204 2492
rect -140 1468 -120 2492
rect 608 2441 712 2839
rect 1388 2788 1408 3812
rect 1472 2788 1492 3812
rect 2220 3761 2324 4159
rect 3000 4108 3020 5132
rect 3084 4108 3104 5132
rect 3832 5081 3936 5280
rect 4612 5132 4716 5280
rect 3423 5080 4345 5081
rect 3423 4160 3424 5080
rect 4344 4160 4345 5080
rect 3423 4159 4345 4160
rect 3000 3812 3104 4108
rect 1811 3760 2733 3761
rect 1811 2840 1812 3760
rect 2732 2840 2733 3760
rect 1811 2839 2733 2840
rect 1388 2492 1492 2788
rect 199 2440 1121 2441
rect 199 1520 200 2440
rect 1120 1520 1121 2440
rect 199 1519 1121 1520
rect -224 1172 -120 1468
rect -1413 1120 -491 1121
rect -1413 200 -1412 1120
rect -492 200 -491 1120
rect -1413 199 -491 200
rect -1836 -148 -1732 148
rect -3025 -200 -2103 -199
rect -3025 -1120 -3024 -200
rect -2104 -1120 -2103 -200
rect -3025 -1121 -2103 -1120
rect -3448 -1468 -3344 -1172
rect -4637 -1520 -3715 -1519
rect -4637 -2440 -4636 -1520
rect -3716 -2440 -3715 -1520
rect -4637 -2441 -3715 -2440
rect -5060 -2788 -4956 -2492
rect -6249 -2840 -5327 -2839
rect -6249 -3760 -6248 -2840
rect -5328 -3760 -5327 -2840
rect -6249 -3761 -5327 -3760
rect -6672 -4108 -6568 -3812
rect -7861 -4160 -6939 -4159
rect -7861 -5080 -7860 -4160
rect -6940 -5080 -6939 -4160
rect -7861 -5081 -6939 -5080
rect -8284 -5280 -8180 -5132
rect -7452 -5280 -7348 -5081
rect -6672 -5132 -6652 -4108
rect -6588 -5132 -6568 -4108
rect -5840 -4159 -5736 -3761
rect -5060 -3812 -5040 -2788
rect -4976 -3812 -4956 -2788
rect -4228 -2839 -4124 -2441
rect -3448 -2492 -3428 -1468
rect -3364 -2492 -3344 -1468
rect -2616 -1519 -2512 -1121
rect -1836 -1172 -1816 -148
rect -1752 -1172 -1732 -148
rect -1004 -199 -900 199
rect -224 148 -204 1172
rect -140 148 -120 1172
rect 608 1121 712 1519
rect 1388 1468 1408 2492
rect 1472 1468 1492 2492
rect 2220 2441 2324 2839
rect 3000 2788 3020 3812
rect 3084 2788 3104 3812
rect 3832 3761 3936 4159
rect 4612 4108 4632 5132
rect 4696 4108 4716 5132
rect 5444 5081 5548 5280
rect 6224 5132 6328 5280
rect 5035 5080 5957 5081
rect 5035 4160 5036 5080
rect 5956 4160 5957 5080
rect 5035 4159 5957 4160
rect 4612 3812 4716 4108
rect 3423 3760 4345 3761
rect 3423 2840 3424 3760
rect 4344 2840 4345 3760
rect 3423 2839 4345 2840
rect 3000 2492 3104 2788
rect 1811 2440 2733 2441
rect 1811 1520 1812 2440
rect 2732 1520 2733 2440
rect 1811 1519 2733 1520
rect 1388 1172 1492 1468
rect 199 1120 1121 1121
rect 199 200 200 1120
rect 1120 200 1121 1120
rect 199 199 1121 200
rect -224 -148 -120 148
rect -1413 -200 -491 -199
rect -1413 -1120 -1412 -200
rect -492 -1120 -491 -200
rect -1413 -1121 -491 -1120
rect -1836 -1468 -1732 -1172
rect -3025 -1520 -2103 -1519
rect -3025 -2440 -3024 -1520
rect -2104 -2440 -2103 -1520
rect -3025 -2441 -2103 -2440
rect -3448 -2788 -3344 -2492
rect -4637 -2840 -3715 -2839
rect -4637 -3760 -4636 -2840
rect -3716 -3760 -3715 -2840
rect -4637 -3761 -3715 -3760
rect -5060 -4108 -4956 -3812
rect -6249 -4160 -5327 -4159
rect -6249 -5080 -6248 -4160
rect -5328 -5080 -5327 -4160
rect -6249 -5081 -5327 -5080
rect -6672 -5280 -6568 -5132
rect -5840 -5280 -5736 -5081
rect -5060 -5132 -5040 -4108
rect -4976 -5132 -4956 -4108
rect -4228 -4159 -4124 -3761
rect -3448 -3812 -3428 -2788
rect -3364 -3812 -3344 -2788
rect -2616 -2839 -2512 -2441
rect -1836 -2492 -1816 -1468
rect -1752 -2492 -1732 -1468
rect -1004 -1519 -900 -1121
rect -224 -1172 -204 -148
rect -140 -1172 -120 -148
rect 608 -199 712 199
rect 1388 148 1408 1172
rect 1472 148 1492 1172
rect 2220 1121 2324 1519
rect 3000 1468 3020 2492
rect 3084 1468 3104 2492
rect 3832 2441 3936 2839
rect 4612 2788 4632 3812
rect 4696 2788 4716 3812
rect 5444 3761 5548 4159
rect 6224 4108 6244 5132
rect 6308 4108 6328 5132
rect 7056 5081 7160 5280
rect 7836 5132 7940 5280
rect 6647 5080 7569 5081
rect 6647 4160 6648 5080
rect 7568 4160 7569 5080
rect 6647 4159 7569 4160
rect 6224 3812 6328 4108
rect 5035 3760 5957 3761
rect 5035 2840 5036 3760
rect 5956 2840 5957 3760
rect 5035 2839 5957 2840
rect 4612 2492 4716 2788
rect 3423 2440 4345 2441
rect 3423 1520 3424 2440
rect 4344 1520 4345 2440
rect 3423 1519 4345 1520
rect 3000 1172 3104 1468
rect 1811 1120 2733 1121
rect 1811 200 1812 1120
rect 2732 200 2733 1120
rect 1811 199 2733 200
rect 1388 -148 1492 148
rect 199 -200 1121 -199
rect 199 -1120 200 -200
rect 1120 -1120 1121 -200
rect 199 -1121 1121 -1120
rect -224 -1468 -120 -1172
rect -1413 -1520 -491 -1519
rect -1413 -2440 -1412 -1520
rect -492 -2440 -491 -1520
rect -1413 -2441 -491 -2440
rect -1836 -2788 -1732 -2492
rect -3025 -2840 -2103 -2839
rect -3025 -3760 -3024 -2840
rect -2104 -3760 -2103 -2840
rect -3025 -3761 -2103 -3760
rect -3448 -4108 -3344 -3812
rect -4637 -4160 -3715 -4159
rect -4637 -5080 -4636 -4160
rect -3716 -5080 -3715 -4160
rect -4637 -5081 -3715 -5080
rect -5060 -5280 -4956 -5132
rect -4228 -5280 -4124 -5081
rect -3448 -5132 -3428 -4108
rect -3364 -5132 -3344 -4108
rect -2616 -4159 -2512 -3761
rect -1836 -3812 -1816 -2788
rect -1752 -3812 -1732 -2788
rect -1004 -2839 -900 -2441
rect -224 -2492 -204 -1468
rect -140 -2492 -120 -1468
rect 608 -1519 712 -1121
rect 1388 -1172 1408 -148
rect 1472 -1172 1492 -148
rect 2220 -199 2324 199
rect 3000 148 3020 1172
rect 3084 148 3104 1172
rect 3832 1121 3936 1519
rect 4612 1468 4632 2492
rect 4696 1468 4716 2492
rect 5444 2441 5548 2839
rect 6224 2788 6244 3812
rect 6308 2788 6328 3812
rect 7056 3761 7160 4159
rect 7836 4108 7856 5132
rect 7920 4108 7940 5132
rect 8668 5081 8772 5280
rect 9448 5132 9552 5280
rect 8259 5080 9181 5081
rect 8259 4160 8260 5080
rect 9180 4160 9181 5080
rect 8259 4159 9181 4160
rect 7836 3812 7940 4108
rect 6647 3760 7569 3761
rect 6647 2840 6648 3760
rect 7568 2840 7569 3760
rect 6647 2839 7569 2840
rect 6224 2492 6328 2788
rect 5035 2440 5957 2441
rect 5035 1520 5036 2440
rect 5956 1520 5957 2440
rect 5035 1519 5957 1520
rect 4612 1172 4716 1468
rect 3423 1120 4345 1121
rect 3423 200 3424 1120
rect 4344 200 4345 1120
rect 3423 199 4345 200
rect 3000 -148 3104 148
rect 1811 -200 2733 -199
rect 1811 -1120 1812 -200
rect 2732 -1120 2733 -200
rect 1811 -1121 2733 -1120
rect 1388 -1468 1492 -1172
rect 199 -1520 1121 -1519
rect 199 -2440 200 -1520
rect 1120 -2440 1121 -1520
rect 199 -2441 1121 -2440
rect -224 -2788 -120 -2492
rect -1413 -2840 -491 -2839
rect -1413 -3760 -1412 -2840
rect -492 -3760 -491 -2840
rect -1413 -3761 -491 -3760
rect -1836 -4108 -1732 -3812
rect -3025 -4160 -2103 -4159
rect -3025 -5080 -3024 -4160
rect -2104 -5080 -2103 -4160
rect -3025 -5081 -2103 -5080
rect -3448 -5280 -3344 -5132
rect -2616 -5280 -2512 -5081
rect -1836 -5132 -1816 -4108
rect -1752 -5132 -1732 -4108
rect -1004 -4159 -900 -3761
rect -224 -3812 -204 -2788
rect -140 -3812 -120 -2788
rect 608 -2839 712 -2441
rect 1388 -2492 1408 -1468
rect 1472 -2492 1492 -1468
rect 2220 -1519 2324 -1121
rect 3000 -1172 3020 -148
rect 3084 -1172 3104 -148
rect 3832 -199 3936 199
rect 4612 148 4632 1172
rect 4696 148 4716 1172
rect 5444 1121 5548 1519
rect 6224 1468 6244 2492
rect 6308 1468 6328 2492
rect 7056 2441 7160 2839
rect 7836 2788 7856 3812
rect 7920 2788 7940 3812
rect 8668 3761 8772 4159
rect 9448 4108 9468 5132
rect 9532 4108 9552 5132
rect 10280 5081 10384 5280
rect 11060 5132 11164 5280
rect 9871 5080 10793 5081
rect 9871 4160 9872 5080
rect 10792 4160 10793 5080
rect 9871 4159 10793 4160
rect 9448 3812 9552 4108
rect 8259 3760 9181 3761
rect 8259 2840 8260 3760
rect 9180 2840 9181 3760
rect 8259 2839 9181 2840
rect 7836 2492 7940 2788
rect 6647 2440 7569 2441
rect 6647 1520 6648 2440
rect 7568 1520 7569 2440
rect 6647 1519 7569 1520
rect 6224 1172 6328 1468
rect 5035 1120 5957 1121
rect 5035 200 5036 1120
rect 5956 200 5957 1120
rect 5035 199 5957 200
rect 4612 -148 4716 148
rect 3423 -200 4345 -199
rect 3423 -1120 3424 -200
rect 4344 -1120 4345 -200
rect 3423 -1121 4345 -1120
rect 3000 -1468 3104 -1172
rect 1811 -1520 2733 -1519
rect 1811 -2440 1812 -1520
rect 2732 -2440 2733 -1520
rect 1811 -2441 2733 -2440
rect 1388 -2788 1492 -2492
rect 199 -2840 1121 -2839
rect 199 -3760 200 -2840
rect 1120 -3760 1121 -2840
rect 199 -3761 1121 -3760
rect -224 -4108 -120 -3812
rect -1413 -4160 -491 -4159
rect -1413 -5080 -1412 -4160
rect -492 -5080 -491 -4160
rect -1413 -5081 -491 -5080
rect -1836 -5280 -1732 -5132
rect -1004 -5280 -900 -5081
rect -224 -5132 -204 -4108
rect -140 -5132 -120 -4108
rect 608 -4159 712 -3761
rect 1388 -3812 1408 -2788
rect 1472 -3812 1492 -2788
rect 2220 -2839 2324 -2441
rect 3000 -2492 3020 -1468
rect 3084 -2492 3104 -1468
rect 3832 -1519 3936 -1121
rect 4612 -1172 4632 -148
rect 4696 -1172 4716 -148
rect 5444 -199 5548 199
rect 6224 148 6244 1172
rect 6308 148 6328 1172
rect 7056 1121 7160 1519
rect 7836 1468 7856 2492
rect 7920 1468 7940 2492
rect 8668 2441 8772 2839
rect 9448 2788 9468 3812
rect 9532 2788 9552 3812
rect 10280 3761 10384 4159
rect 11060 4108 11080 5132
rect 11144 4108 11164 5132
rect 11892 5081 11996 5280
rect 12672 5132 12776 5280
rect 11483 5080 12405 5081
rect 11483 4160 11484 5080
rect 12404 4160 12405 5080
rect 11483 4159 12405 4160
rect 11060 3812 11164 4108
rect 9871 3760 10793 3761
rect 9871 2840 9872 3760
rect 10792 2840 10793 3760
rect 9871 2839 10793 2840
rect 9448 2492 9552 2788
rect 8259 2440 9181 2441
rect 8259 1520 8260 2440
rect 9180 1520 9181 2440
rect 8259 1519 9181 1520
rect 7836 1172 7940 1468
rect 6647 1120 7569 1121
rect 6647 200 6648 1120
rect 7568 200 7569 1120
rect 6647 199 7569 200
rect 6224 -148 6328 148
rect 5035 -200 5957 -199
rect 5035 -1120 5036 -200
rect 5956 -1120 5957 -200
rect 5035 -1121 5957 -1120
rect 4612 -1468 4716 -1172
rect 3423 -1520 4345 -1519
rect 3423 -2440 3424 -1520
rect 4344 -2440 4345 -1520
rect 3423 -2441 4345 -2440
rect 3000 -2788 3104 -2492
rect 1811 -2840 2733 -2839
rect 1811 -3760 1812 -2840
rect 2732 -3760 2733 -2840
rect 1811 -3761 2733 -3760
rect 1388 -4108 1492 -3812
rect 199 -4160 1121 -4159
rect 199 -5080 200 -4160
rect 1120 -5080 1121 -4160
rect 199 -5081 1121 -5080
rect -224 -5280 -120 -5132
rect 608 -5280 712 -5081
rect 1388 -5132 1408 -4108
rect 1472 -5132 1492 -4108
rect 2220 -4159 2324 -3761
rect 3000 -3812 3020 -2788
rect 3084 -3812 3104 -2788
rect 3832 -2839 3936 -2441
rect 4612 -2492 4632 -1468
rect 4696 -2492 4716 -1468
rect 5444 -1519 5548 -1121
rect 6224 -1172 6244 -148
rect 6308 -1172 6328 -148
rect 7056 -199 7160 199
rect 7836 148 7856 1172
rect 7920 148 7940 1172
rect 8668 1121 8772 1519
rect 9448 1468 9468 2492
rect 9532 1468 9552 2492
rect 10280 2441 10384 2839
rect 11060 2788 11080 3812
rect 11144 2788 11164 3812
rect 11892 3761 11996 4159
rect 12672 4108 12692 5132
rect 12756 4108 12776 5132
rect 12672 3812 12776 4108
rect 11483 3760 12405 3761
rect 11483 2840 11484 3760
rect 12404 2840 12405 3760
rect 11483 2839 12405 2840
rect 11060 2492 11164 2788
rect 9871 2440 10793 2441
rect 9871 1520 9872 2440
rect 10792 1520 10793 2440
rect 9871 1519 10793 1520
rect 9448 1172 9552 1468
rect 8259 1120 9181 1121
rect 8259 200 8260 1120
rect 9180 200 9181 1120
rect 8259 199 9181 200
rect 7836 -148 7940 148
rect 6647 -200 7569 -199
rect 6647 -1120 6648 -200
rect 7568 -1120 7569 -200
rect 6647 -1121 7569 -1120
rect 6224 -1468 6328 -1172
rect 5035 -1520 5957 -1519
rect 5035 -2440 5036 -1520
rect 5956 -2440 5957 -1520
rect 5035 -2441 5957 -2440
rect 4612 -2788 4716 -2492
rect 3423 -2840 4345 -2839
rect 3423 -3760 3424 -2840
rect 4344 -3760 4345 -2840
rect 3423 -3761 4345 -3760
rect 3000 -4108 3104 -3812
rect 1811 -4160 2733 -4159
rect 1811 -5080 1812 -4160
rect 2732 -5080 2733 -4160
rect 1811 -5081 2733 -5080
rect 1388 -5280 1492 -5132
rect 2220 -5280 2324 -5081
rect 3000 -5132 3020 -4108
rect 3084 -5132 3104 -4108
rect 3832 -4159 3936 -3761
rect 4612 -3812 4632 -2788
rect 4696 -3812 4716 -2788
rect 5444 -2839 5548 -2441
rect 6224 -2492 6244 -1468
rect 6308 -2492 6328 -1468
rect 7056 -1519 7160 -1121
rect 7836 -1172 7856 -148
rect 7920 -1172 7940 -148
rect 8668 -199 8772 199
rect 9448 148 9468 1172
rect 9532 148 9552 1172
rect 10280 1121 10384 1519
rect 11060 1468 11080 2492
rect 11144 1468 11164 2492
rect 11892 2441 11996 2839
rect 12672 2788 12692 3812
rect 12756 2788 12776 3812
rect 12672 2492 12776 2788
rect 11483 2440 12405 2441
rect 11483 1520 11484 2440
rect 12404 1520 12405 2440
rect 11483 1519 12405 1520
rect 11060 1172 11164 1468
rect 9871 1120 10793 1121
rect 9871 200 9872 1120
rect 10792 200 10793 1120
rect 9871 199 10793 200
rect 9448 -148 9552 148
rect 8259 -200 9181 -199
rect 8259 -1120 8260 -200
rect 9180 -1120 9181 -200
rect 8259 -1121 9181 -1120
rect 7836 -1468 7940 -1172
rect 6647 -1520 7569 -1519
rect 6647 -2440 6648 -1520
rect 7568 -2440 7569 -1520
rect 6647 -2441 7569 -2440
rect 6224 -2788 6328 -2492
rect 5035 -2840 5957 -2839
rect 5035 -3760 5036 -2840
rect 5956 -3760 5957 -2840
rect 5035 -3761 5957 -3760
rect 4612 -4108 4716 -3812
rect 3423 -4160 4345 -4159
rect 3423 -5080 3424 -4160
rect 4344 -5080 4345 -4160
rect 3423 -5081 4345 -5080
rect 3000 -5280 3104 -5132
rect 3832 -5280 3936 -5081
rect 4612 -5132 4632 -4108
rect 4696 -5132 4716 -4108
rect 5444 -4159 5548 -3761
rect 6224 -3812 6244 -2788
rect 6308 -3812 6328 -2788
rect 7056 -2839 7160 -2441
rect 7836 -2492 7856 -1468
rect 7920 -2492 7940 -1468
rect 8668 -1519 8772 -1121
rect 9448 -1172 9468 -148
rect 9532 -1172 9552 -148
rect 10280 -199 10384 199
rect 11060 148 11080 1172
rect 11144 148 11164 1172
rect 11892 1121 11996 1519
rect 12672 1468 12692 2492
rect 12756 1468 12776 2492
rect 12672 1172 12776 1468
rect 11483 1120 12405 1121
rect 11483 200 11484 1120
rect 12404 200 12405 1120
rect 11483 199 12405 200
rect 11060 -148 11164 148
rect 9871 -200 10793 -199
rect 9871 -1120 9872 -200
rect 10792 -1120 10793 -200
rect 9871 -1121 10793 -1120
rect 9448 -1468 9552 -1172
rect 8259 -1520 9181 -1519
rect 8259 -2440 8260 -1520
rect 9180 -2440 9181 -1520
rect 8259 -2441 9181 -2440
rect 7836 -2788 7940 -2492
rect 6647 -2840 7569 -2839
rect 6647 -3760 6648 -2840
rect 7568 -3760 7569 -2840
rect 6647 -3761 7569 -3760
rect 6224 -4108 6328 -3812
rect 5035 -4160 5957 -4159
rect 5035 -5080 5036 -4160
rect 5956 -5080 5957 -4160
rect 5035 -5081 5957 -5080
rect 4612 -5280 4716 -5132
rect 5444 -5280 5548 -5081
rect 6224 -5132 6244 -4108
rect 6308 -5132 6328 -4108
rect 7056 -4159 7160 -3761
rect 7836 -3812 7856 -2788
rect 7920 -3812 7940 -2788
rect 8668 -2839 8772 -2441
rect 9448 -2492 9468 -1468
rect 9532 -2492 9552 -1468
rect 10280 -1519 10384 -1121
rect 11060 -1172 11080 -148
rect 11144 -1172 11164 -148
rect 11892 -199 11996 199
rect 12672 148 12692 1172
rect 12756 148 12776 1172
rect 12672 -148 12776 148
rect 11483 -200 12405 -199
rect 11483 -1120 11484 -200
rect 12404 -1120 12405 -200
rect 11483 -1121 12405 -1120
rect 11060 -1468 11164 -1172
rect 9871 -1520 10793 -1519
rect 9871 -2440 9872 -1520
rect 10792 -2440 10793 -1520
rect 9871 -2441 10793 -2440
rect 9448 -2788 9552 -2492
rect 8259 -2840 9181 -2839
rect 8259 -3760 8260 -2840
rect 9180 -3760 9181 -2840
rect 8259 -3761 9181 -3760
rect 7836 -4108 7940 -3812
rect 6647 -4160 7569 -4159
rect 6647 -5080 6648 -4160
rect 7568 -5080 7569 -4160
rect 6647 -5081 7569 -5080
rect 6224 -5280 6328 -5132
rect 7056 -5280 7160 -5081
rect 7836 -5132 7856 -4108
rect 7920 -5132 7940 -4108
rect 8668 -4159 8772 -3761
rect 9448 -3812 9468 -2788
rect 9532 -3812 9552 -2788
rect 10280 -2839 10384 -2441
rect 11060 -2492 11080 -1468
rect 11144 -2492 11164 -1468
rect 11892 -1519 11996 -1121
rect 12672 -1172 12692 -148
rect 12756 -1172 12776 -148
rect 12672 -1468 12776 -1172
rect 11483 -1520 12405 -1519
rect 11483 -2440 11484 -1520
rect 12404 -2440 12405 -1520
rect 11483 -2441 12405 -2440
rect 11060 -2788 11164 -2492
rect 9871 -2840 10793 -2839
rect 9871 -3760 9872 -2840
rect 10792 -3760 10793 -2840
rect 9871 -3761 10793 -3760
rect 9448 -4108 9552 -3812
rect 8259 -4160 9181 -4159
rect 8259 -5080 8260 -4160
rect 9180 -5080 9181 -4160
rect 8259 -5081 9181 -5080
rect 7836 -5280 7940 -5132
rect 8668 -5280 8772 -5081
rect 9448 -5132 9468 -4108
rect 9532 -5132 9552 -4108
rect 10280 -4159 10384 -3761
rect 11060 -3812 11080 -2788
rect 11144 -3812 11164 -2788
rect 11892 -2839 11996 -2441
rect 12672 -2492 12692 -1468
rect 12756 -2492 12776 -1468
rect 12672 -2788 12776 -2492
rect 11483 -2840 12405 -2839
rect 11483 -3760 11484 -2840
rect 12404 -3760 12405 -2840
rect 11483 -3761 12405 -3760
rect 11060 -4108 11164 -3812
rect 9871 -4160 10793 -4159
rect 9871 -5080 9872 -4160
rect 10792 -5080 10793 -4160
rect 9871 -5081 10793 -5080
rect 9448 -5280 9552 -5132
rect 10280 -5280 10384 -5081
rect 11060 -5132 11080 -4108
rect 11144 -5132 11164 -4108
rect 11892 -4159 11996 -3761
rect 12672 -3812 12692 -2788
rect 12756 -3812 12776 -2788
rect 12672 -4108 12776 -3812
rect 11483 -4160 12405 -4159
rect 11483 -5080 11484 -4160
rect 12404 -5080 12405 -4160
rect 11483 -5081 12405 -5080
rect 11060 -5280 11164 -5132
rect 11892 -5280 11996 -5081
rect 12672 -5132 12692 -4108
rect 12756 -5132 12776 -4108
rect 12672 -5280 12776 -5132
<< properties >>
string FIXED_BBOX 11404 4080 12484 5160
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5.0 l 5.0 val 53.8 carea 2.00 cperi 0.19 nx 16 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

** sch_path: /home/ttuser/Documents/SARADC/xschem/cap128/cap128.sch
**.subckt cap128 bottom top
*.ipin bottom
*.ipin top
XC12 top bottom sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=128 m=128
**.ends
.end

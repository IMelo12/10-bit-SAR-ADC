** sch_path: /home/ttuser/Documents/SARADC/xschem/cap4/cap4.sch
**.subckt cap4 bottom top
*.ipin bottom
*.ipin top
XC12 top bottom sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=4 m=4
**.ends
.end

magic
tech sky130A
magscale 1 2
timestamp 1754941660
<< metal3 >>
rect -686 5132 686 5160
rect -686 4108 602 5132
rect 666 4108 686 5132
rect -686 4080 686 4108
rect -686 3812 686 3840
rect -686 2788 602 3812
rect 666 2788 686 3812
rect -686 2760 686 2788
rect -686 2492 686 2520
rect -686 1468 602 2492
rect 666 1468 686 2492
rect -686 1440 686 1468
rect -686 1172 686 1200
rect -686 148 602 1172
rect 666 148 686 1172
rect -686 120 686 148
rect -686 -148 686 -120
rect -686 -1172 602 -148
rect 666 -1172 686 -148
rect -686 -1200 686 -1172
rect -686 -1468 686 -1440
rect -686 -2492 602 -1468
rect 666 -2492 686 -1468
rect -686 -2520 686 -2492
rect -686 -2788 686 -2760
rect -686 -3812 602 -2788
rect 666 -3812 686 -2788
rect -686 -3840 686 -3812
rect -686 -4108 686 -4080
rect -686 -5132 602 -4108
rect 666 -5132 686 -4108
rect -686 -5160 686 -5132
<< via3 >>
rect 602 4108 666 5132
rect 602 2788 666 3812
rect 602 1468 666 2492
rect 602 148 666 1172
rect 602 -1172 666 -148
rect 602 -2492 666 -1468
rect 602 -3812 666 -2788
rect 602 -5132 666 -4108
<< mimcap >>
rect -646 5080 354 5120
rect -646 4160 -606 5080
rect 314 4160 354 5080
rect -646 4120 354 4160
rect -646 3760 354 3800
rect -646 2840 -606 3760
rect 314 2840 354 3760
rect -646 2800 354 2840
rect -646 2440 354 2480
rect -646 1520 -606 2440
rect 314 1520 354 2440
rect -646 1480 354 1520
rect -646 1120 354 1160
rect -646 200 -606 1120
rect 314 200 354 1120
rect -646 160 354 200
rect -646 -200 354 -160
rect -646 -1120 -606 -200
rect 314 -1120 354 -200
rect -646 -1160 354 -1120
rect -646 -1520 354 -1480
rect -646 -2440 -606 -1520
rect 314 -2440 354 -1520
rect -646 -2480 354 -2440
rect -646 -2840 354 -2800
rect -646 -3760 -606 -2840
rect 314 -3760 354 -2840
rect -646 -3800 354 -3760
rect -646 -4160 354 -4120
rect -646 -5080 -606 -4160
rect 314 -5080 354 -4160
rect -646 -5120 354 -5080
<< mimcapcontact >>
rect -606 4160 314 5080
rect -606 2840 314 3760
rect -606 1520 314 2440
rect -606 200 314 1120
rect -606 -1120 314 -200
rect -606 -2440 314 -1520
rect -606 -3760 314 -2840
rect -606 -5080 314 -4160
<< metal4 >>
rect -198 5081 -94 5280
rect 582 5132 686 5280
rect -607 5080 315 5081
rect -607 4160 -606 5080
rect 314 4160 315 5080
rect -607 4159 315 4160
rect -198 3761 -94 4159
rect 582 4108 602 5132
rect 666 4108 686 5132
rect 582 3812 686 4108
rect -607 3760 315 3761
rect -607 2840 -606 3760
rect 314 2840 315 3760
rect -607 2839 315 2840
rect -198 2441 -94 2839
rect 582 2788 602 3812
rect 666 2788 686 3812
rect 582 2492 686 2788
rect -607 2440 315 2441
rect -607 1520 -606 2440
rect 314 1520 315 2440
rect -607 1519 315 1520
rect -198 1121 -94 1519
rect 582 1468 602 2492
rect 666 1468 686 2492
rect 582 1172 686 1468
rect -607 1120 315 1121
rect -607 200 -606 1120
rect 314 200 315 1120
rect -607 199 315 200
rect -198 -199 -94 199
rect 582 148 602 1172
rect 666 148 686 1172
rect 582 -148 686 148
rect -607 -200 315 -199
rect -607 -1120 -606 -200
rect 314 -1120 315 -200
rect -607 -1121 315 -1120
rect -198 -1519 -94 -1121
rect 582 -1172 602 -148
rect 666 -1172 686 -148
rect 582 -1468 686 -1172
rect -607 -1520 315 -1519
rect -607 -2440 -606 -1520
rect 314 -2440 315 -1520
rect -607 -2441 315 -2440
rect -198 -2839 -94 -2441
rect 582 -2492 602 -1468
rect 666 -2492 686 -1468
rect 582 -2788 686 -2492
rect -607 -2840 315 -2839
rect -607 -3760 -606 -2840
rect 314 -3760 315 -2840
rect -607 -3761 315 -3760
rect -198 -4159 -94 -3761
rect 582 -3812 602 -2788
rect 666 -3812 686 -2788
rect 582 -4108 686 -3812
rect -607 -4160 315 -4159
rect -607 -5080 -606 -4160
rect 314 -5080 315 -4160
rect -607 -5081 315 -5080
rect -198 -5280 -94 -5081
rect 582 -5132 602 -4108
rect 666 -5132 686 -4108
rect 582 -5280 686 -5132
<< properties >>
string FIXED_BBOX -686 4080 394 5160
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5.0 l 5.0 val 53.8 carea 2.00 cperi 0.19 nx 1 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

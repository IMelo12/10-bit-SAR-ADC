** sch_path: /home/ttuser/Documents/SARADC/xschem/cap8/cap8.sch
**.subckt cap8 bottom top
*.ipin bottom
*.ipin top
XC12 top bottom sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=8 m=8
**.ends
.end

** sch_path: /home/ttuser/Documents/SARADC/xschem/cap32/cap32.sch
**.subckt cap32 bottom top
*.ipin bottom
*.ipin top
XC12 top bottom sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=32 m=32
**.ends
.end

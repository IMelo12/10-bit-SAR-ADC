magic
tech sky130A
magscale 1 2
timestamp 1754899758
<< metal3 >>
rect -12776 1172 -11404 1200
rect -12776 148 -11488 1172
rect -11424 148 -11404 1172
rect -12776 120 -11404 148
rect -11164 1172 -9792 1200
rect -11164 148 -9876 1172
rect -9812 148 -9792 1172
rect -11164 120 -9792 148
rect -9552 1172 -8180 1200
rect -9552 148 -8264 1172
rect -8200 148 -8180 1172
rect -9552 120 -8180 148
rect -7940 1172 -6568 1200
rect -7940 148 -6652 1172
rect -6588 148 -6568 1172
rect -7940 120 -6568 148
rect -6328 1172 -4956 1200
rect -6328 148 -5040 1172
rect -4976 148 -4956 1172
rect -6328 120 -4956 148
rect -4716 1172 -3344 1200
rect -4716 148 -3428 1172
rect -3364 148 -3344 1172
rect -4716 120 -3344 148
rect -3104 1172 -1732 1200
rect -3104 148 -1816 1172
rect -1752 148 -1732 1172
rect -3104 120 -1732 148
rect -1492 1172 -120 1200
rect -1492 148 -204 1172
rect -140 148 -120 1172
rect -1492 120 -120 148
rect 120 1172 1492 1200
rect 120 148 1408 1172
rect 1472 148 1492 1172
rect 120 120 1492 148
rect 1732 1172 3104 1200
rect 1732 148 3020 1172
rect 3084 148 3104 1172
rect 1732 120 3104 148
rect 3344 1172 4716 1200
rect 3344 148 4632 1172
rect 4696 148 4716 1172
rect 3344 120 4716 148
rect 4956 1172 6328 1200
rect 4956 148 6244 1172
rect 6308 148 6328 1172
rect 4956 120 6328 148
rect 6568 1172 7940 1200
rect 6568 148 7856 1172
rect 7920 148 7940 1172
rect 6568 120 7940 148
rect 8180 1172 9552 1200
rect 8180 148 9468 1172
rect 9532 148 9552 1172
rect 8180 120 9552 148
rect 9792 1172 11164 1200
rect 9792 148 11080 1172
rect 11144 148 11164 1172
rect 9792 120 11164 148
rect 11404 1172 12776 1200
rect 11404 148 12692 1172
rect 12756 148 12776 1172
rect 11404 120 12776 148
rect -12776 -148 -11404 -120
rect -12776 -1172 -11488 -148
rect -11424 -1172 -11404 -148
rect -12776 -1200 -11404 -1172
rect -11164 -148 -9792 -120
rect -11164 -1172 -9876 -148
rect -9812 -1172 -9792 -148
rect -11164 -1200 -9792 -1172
rect -9552 -148 -8180 -120
rect -9552 -1172 -8264 -148
rect -8200 -1172 -8180 -148
rect -9552 -1200 -8180 -1172
rect -7940 -148 -6568 -120
rect -7940 -1172 -6652 -148
rect -6588 -1172 -6568 -148
rect -7940 -1200 -6568 -1172
rect -6328 -148 -4956 -120
rect -6328 -1172 -5040 -148
rect -4976 -1172 -4956 -148
rect -6328 -1200 -4956 -1172
rect -4716 -148 -3344 -120
rect -4716 -1172 -3428 -148
rect -3364 -1172 -3344 -148
rect -4716 -1200 -3344 -1172
rect -3104 -148 -1732 -120
rect -3104 -1172 -1816 -148
rect -1752 -1172 -1732 -148
rect -3104 -1200 -1732 -1172
rect -1492 -148 -120 -120
rect -1492 -1172 -204 -148
rect -140 -1172 -120 -148
rect -1492 -1200 -120 -1172
rect 120 -148 1492 -120
rect 120 -1172 1408 -148
rect 1472 -1172 1492 -148
rect 120 -1200 1492 -1172
rect 1732 -148 3104 -120
rect 1732 -1172 3020 -148
rect 3084 -1172 3104 -148
rect 1732 -1200 3104 -1172
rect 3344 -148 4716 -120
rect 3344 -1172 4632 -148
rect 4696 -1172 4716 -148
rect 3344 -1200 4716 -1172
rect 4956 -148 6328 -120
rect 4956 -1172 6244 -148
rect 6308 -1172 6328 -148
rect 4956 -1200 6328 -1172
rect 6568 -148 7940 -120
rect 6568 -1172 7856 -148
rect 7920 -1172 7940 -148
rect 6568 -1200 7940 -1172
rect 8180 -148 9552 -120
rect 8180 -1172 9468 -148
rect 9532 -1172 9552 -148
rect 8180 -1200 9552 -1172
rect 9792 -148 11164 -120
rect 9792 -1172 11080 -148
rect 11144 -1172 11164 -148
rect 9792 -1200 11164 -1172
rect 11404 -148 12776 -120
rect 11404 -1172 12692 -148
rect 12756 -1172 12776 -148
rect 11404 -1200 12776 -1172
<< via3 >>
rect -11488 148 -11424 1172
rect -9876 148 -9812 1172
rect -8264 148 -8200 1172
rect -6652 148 -6588 1172
rect -5040 148 -4976 1172
rect -3428 148 -3364 1172
rect -1816 148 -1752 1172
rect -204 148 -140 1172
rect 1408 148 1472 1172
rect 3020 148 3084 1172
rect 4632 148 4696 1172
rect 6244 148 6308 1172
rect 7856 148 7920 1172
rect 9468 148 9532 1172
rect 11080 148 11144 1172
rect 12692 148 12756 1172
rect -11488 -1172 -11424 -148
rect -9876 -1172 -9812 -148
rect -8264 -1172 -8200 -148
rect -6652 -1172 -6588 -148
rect -5040 -1172 -4976 -148
rect -3428 -1172 -3364 -148
rect -1816 -1172 -1752 -148
rect -204 -1172 -140 -148
rect 1408 -1172 1472 -148
rect 3020 -1172 3084 -148
rect 4632 -1172 4696 -148
rect 6244 -1172 6308 -148
rect 7856 -1172 7920 -148
rect 9468 -1172 9532 -148
rect 11080 -1172 11144 -148
rect 12692 -1172 12756 -148
<< mimcap >>
rect -12736 1120 -11736 1160
rect -12736 200 -12696 1120
rect -11776 200 -11736 1120
rect -12736 160 -11736 200
rect -11124 1120 -10124 1160
rect -11124 200 -11084 1120
rect -10164 200 -10124 1120
rect -11124 160 -10124 200
rect -9512 1120 -8512 1160
rect -9512 200 -9472 1120
rect -8552 200 -8512 1120
rect -9512 160 -8512 200
rect -7900 1120 -6900 1160
rect -7900 200 -7860 1120
rect -6940 200 -6900 1120
rect -7900 160 -6900 200
rect -6288 1120 -5288 1160
rect -6288 200 -6248 1120
rect -5328 200 -5288 1120
rect -6288 160 -5288 200
rect -4676 1120 -3676 1160
rect -4676 200 -4636 1120
rect -3716 200 -3676 1120
rect -4676 160 -3676 200
rect -3064 1120 -2064 1160
rect -3064 200 -3024 1120
rect -2104 200 -2064 1120
rect -3064 160 -2064 200
rect -1452 1120 -452 1160
rect -1452 200 -1412 1120
rect -492 200 -452 1120
rect -1452 160 -452 200
rect 160 1120 1160 1160
rect 160 200 200 1120
rect 1120 200 1160 1120
rect 160 160 1160 200
rect 1772 1120 2772 1160
rect 1772 200 1812 1120
rect 2732 200 2772 1120
rect 1772 160 2772 200
rect 3384 1120 4384 1160
rect 3384 200 3424 1120
rect 4344 200 4384 1120
rect 3384 160 4384 200
rect 4996 1120 5996 1160
rect 4996 200 5036 1120
rect 5956 200 5996 1120
rect 4996 160 5996 200
rect 6608 1120 7608 1160
rect 6608 200 6648 1120
rect 7568 200 7608 1120
rect 6608 160 7608 200
rect 8220 1120 9220 1160
rect 8220 200 8260 1120
rect 9180 200 9220 1120
rect 8220 160 9220 200
rect 9832 1120 10832 1160
rect 9832 200 9872 1120
rect 10792 200 10832 1120
rect 9832 160 10832 200
rect 11444 1120 12444 1160
rect 11444 200 11484 1120
rect 12404 200 12444 1120
rect 11444 160 12444 200
rect -12736 -200 -11736 -160
rect -12736 -1120 -12696 -200
rect -11776 -1120 -11736 -200
rect -12736 -1160 -11736 -1120
rect -11124 -200 -10124 -160
rect -11124 -1120 -11084 -200
rect -10164 -1120 -10124 -200
rect -11124 -1160 -10124 -1120
rect -9512 -200 -8512 -160
rect -9512 -1120 -9472 -200
rect -8552 -1120 -8512 -200
rect -9512 -1160 -8512 -1120
rect -7900 -200 -6900 -160
rect -7900 -1120 -7860 -200
rect -6940 -1120 -6900 -200
rect -7900 -1160 -6900 -1120
rect -6288 -200 -5288 -160
rect -6288 -1120 -6248 -200
rect -5328 -1120 -5288 -200
rect -6288 -1160 -5288 -1120
rect -4676 -200 -3676 -160
rect -4676 -1120 -4636 -200
rect -3716 -1120 -3676 -200
rect -4676 -1160 -3676 -1120
rect -3064 -200 -2064 -160
rect -3064 -1120 -3024 -200
rect -2104 -1120 -2064 -200
rect -3064 -1160 -2064 -1120
rect -1452 -200 -452 -160
rect -1452 -1120 -1412 -200
rect -492 -1120 -452 -200
rect -1452 -1160 -452 -1120
rect 160 -200 1160 -160
rect 160 -1120 200 -200
rect 1120 -1120 1160 -200
rect 160 -1160 1160 -1120
rect 1772 -200 2772 -160
rect 1772 -1120 1812 -200
rect 2732 -1120 2772 -200
rect 1772 -1160 2772 -1120
rect 3384 -200 4384 -160
rect 3384 -1120 3424 -200
rect 4344 -1120 4384 -200
rect 3384 -1160 4384 -1120
rect 4996 -200 5996 -160
rect 4996 -1120 5036 -200
rect 5956 -1120 5996 -200
rect 4996 -1160 5996 -1120
rect 6608 -200 7608 -160
rect 6608 -1120 6648 -200
rect 7568 -1120 7608 -200
rect 6608 -1160 7608 -1120
rect 8220 -200 9220 -160
rect 8220 -1120 8260 -200
rect 9180 -1120 9220 -200
rect 8220 -1160 9220 -1120
rect 9832 -200 10832 -160
rect 9832 -1120 9872 -200
rect 10792 -1120 10832 -200
rect 9832 -1160 10832 -1120
rect 11444 -200 12444 -160
rect 11444 -1120 11484 -200
rect 12404 -1120 12444 -200
rect 11444 -1160 12444 -1120
<< mimcapcontact >>
rect -12696 200 -11776 1120
rect -11084 200 -10164 1120
rect -9472 200 -8552 1120
rect -7860 200 -6940 1120
rect -6248 200 -5328 1120
rect -4636 200 -3716 1120
rect -3024 200 -2104 1120
rect -1412 200 -492 1120
rect 200 200 1120 1120
rect 1812 200 2732 1120
rect 3424 200 4344 1120
rect 5036 200 5956 1120
rect 6648 200 7568 1120
rect 8260 200 9180 1120
rect 9872 200 10792 1120
rect 11484 200 12404 1120
rect -12696 -1120 -11776 -200
rect -11084 -1120 -10164 -200
rect -9472 -1120 -8552 -200
rect -7860 -1120 -6940 -200
rect -6248 -1120 -5328 -200
rect -4636 -1120 -3716 -200
rect -3024 -1120 -2104 -200
rect -1412 -1120 -492 -200
rect 200 -1120 1120 -200
rect 1812 -1120 2732 -200
rect 3424 -1120 4344 -200
rect 5036 -1120 5956 -200
rect 6648 -1120 7568 -200
rect 8260 -1120 9180 -200
rect 9872 -1120 10792 -200
rect 11484 -1120 12404 -200
<< metal4 >>
rect -12288 1121 -12184 1320
rect -11508 1172 -11404 1320
rect -12697 1120 -11775 1121
rect -12697 200 -12696 1120
rect -11776 200 -11775 1120
rect -12697 199 -11775 200
rect -12288 -199 -12184 199
rect -11508 148 -11488 1172
rect -11424 148 -11404 1172
rect -10676 1121 -10572 1320
rect -9896 1172 -9792 1320
rect -11085 1120 -10163 1121
rect -11085 200 -11084 1120
rect -10164 200 -10163 1120
rect -11085 199 -10163 200
rect -11508 -148 -11404 148
rect -12697 -200 -11775 -199
rect -12697 -1120 -12696 -200
rect -11776 -1120 -11775 -200
rect -12697 -1121 -11775 -1120
rect -12288 -1320 -12184 -1121
rect -11508 -1172 -11488 -148
rect -11424 -1172 -11404 -148
rect -10676 -199 -10572 199
rect -9896 148 -9876 1172
rect -9812 148 -9792 1172
rect -9064 1121 -8960 1320
rect -8284 1172 -8180 1320
rect -9473 1120 -8551 1121
rect -9473 200 -9472 1120
rect -8552 200 -8551 1120
rect -9473 199 -8551 200
rect -9896 -148 -9792 148
rect -11085 -200 -10163 -199
rect -11085 -1120 -11084 -200
rect -10164 -1120 -10163 -200
rect -11085 -1121 -10163 -1120
rect -11508 -1320 -11404 -1172
rect -10676 -1320 -10572 -1121
rect -9896 -1172 -9876 -148
rect -9812 -1172 -9792 -148
rect -9064 -199 -8960 199
rect -8284 148 -8264 1172
rect -8200 148 -8180 1172
rect -7452 1121 -7348 1320
rect -6672 1172 -6568 1320
rect -7861 1120 -6939 1121
rect -7861 200 -7860 1120
rect -6940 200 -6939 1120
rect -7861 199 -6939 200
rect -8284 -148 -8180 148
rect -9473 -200 -8551 -199
rect -9473 -1120 -9472 -200
rect -8552 -1120 -8551 -200
rect -9473 -1121 -8551 -1120
rect -9896 -1320 -9792 -1172
rect -9064 -1320 -8960 -1121
rect -8284 -1172 -8264 -148
rect -8200 -1172 -8180 -148
rect -7452 -199 -7348 199
rect -6672 148 -6652 1172
rect -6588 148 -6568 1172
rect -5840 1121 -5736 1320
rect -5060 1172 -4956 1320
rect -6249 1120 -5327 1121
rect -6249 200 -6248 1120
rect -5328 200 -5327 1120
rect -6249 199 -5327 200
rect -6672 -148 -6568 148
rect -7861 -200 -6939 -199
rect -7861 -1120 -7860 -200
rect -6940 -1120 -6939 -200
rect -7861 -1121 -6939 -1120
rect -8284 -1320 -8180 -1172
rect -7452 -1320 -7348 -1121
rect -6672 -1172 -6652 -148
rect -6588 -1172 -6568 -148
rect -5840 -199 -5736 199
rect -5060 148 -5040 1172
rect -4976 148 -4956 1172
rect -4228 1121 -4124 1320
rect -3448 1172 -3344 1320
rect -4637 1120 -3715 1121
rect -4637 200 -4636 1120
rect -3716 200 -3715 1120
rect -4637 199 -3715 200
rect -5060 -148 -4956 148
rect -6249 -200 -5327 -199
rect -6249 -1120 -6248 -200
rect -5328 -1120 -5327 -200
rect -6249 -1121 -5327 -1120
rect -6672 -1320 -6568 -1172
rect -5840 -1320 -5736 -1121
rect -5060 -1172 -5040 -148
rect -4976 -1172 -4956 -148
rect -4228 -199 -4124 199
rect -3448 148 -3428 1172
rect -3364 148 -3344 1172
rect -2616 1121 -2512 1320
rect -1836 1172 -1732 1320
rect -3025 1120 -2103 1121
rect -3025 200 -3024 1120
rect -2104 200 -2103 1120
rect -3025 199 -2103 200
rect -3448 -148 -3344 148
rect -4637 -200 -3715 -199
rect -4637 -1120 -4636 -200
rect -3716 -1120 -3715 -200
rect -4637 -1121 -3715 -1120
rect -5060 -1320 -4956 -1172
rect -4228 -1320 -4124 -1121
rect -3448 -1172 -3428 -148
rect -3364 -1172 -3344 -148
rect -2616 -199 -2512 199
rect -1836 148 -1816 1172
rect -1752 148 -1732 1172
rect -1004 1121 -900 1320
rect -224 1172 -120 1320
rect -1413 1120 -491 1121
rect -1413 200 -1412 1120
rect -492 200 -491 1120
rect -1413 199 -491 200
rect -1836 -148 -1732 148
rect -3025 -200 -2103 -199
rect -3025 -1120 -3024 -200
rect -2104 -1120 -2103 -200
rect -3025 -1121 -2103 -1120
rect -3448 -1320 -3344 -1172
rect -2616 -1320 -2512 -1121
rect -1836 -1172 -1816 -148
rect -1752 -1172 -1732 -148
rect -1004 -199 -900 199
rect -224 148 -204 1172
rect -140 148 -120 1172
rect 608 1121 712 1320
rect 1388 1172 1492 1320
rect 199 1120 1121 1121
rect 199 200 200 1120
rect 1120 200 1121 1120
rect 199 199 1121 200
rect -224 -148 -120 148
rect -1413 -200 -491 -199
rect -1413 -1120 -1412 -200
rect -492 -1120 -491 -200
rect -1413 -1121 -491 -1120
rect -1836 -1320 -1732 -1172
rect -1004 -1320 -900 -1121
rect -224 -1172 -204 -148
rect -140 -1172 -120 -148
rect 608 -199 712 199
rect 1388 148 1408 1172
rect 1472 148 1492 1172
rect 2220 1121 2324 1320
rect 3000 1172 3104 1320
rect 1811 1120 2733 1121
rect 1811 200 1812 1120
rect 2732 200 2733 1120
rect 1811 199 2733 200
rect 1388 -148 1492 148
rect 199 -200 1121 -199
rect 199 -1120 200 -200
rect 1120 -1120 1121 -200
rect 199 -1121 1121 -1120
rect -224 -1320 -120 -1172
rect 608 -1320 712 -1121
rect 1388 -1172 1408 -148
rect 1472 -1172 1492 -148
rect 2220 -199 2324 199
rect 3000 148 3020 1172
rect 3084 148 3104 1172
rect 3832 1121 3936 1320
rect 4612 1172 4716 1320
rect 3423 1120 4345 1121
rect 3423 200 3424 1120
rect 4344 200 4345 1120
rect 3423 199 4345 200
rect 3000 -148 3104 148
rect 1811 -200 2733 -199
rect 1811 -1120 1812 -200
rect 2732 -1120 2733 -200
rect 1811 -1121 2733 -1120
rect 1388 -1320 1492 -1172
rect 2220 -1320 2324 -1121
rect 3000 -1172 3020 -148
rect 3084 -1172 3104 -148
rect 3832 -199 3936 199
rect 4612 148 4632 1172
rect 4696 148 4716 1172
rect 5444 1121 5548 1320
rect 6224 1172 6328 1320
rect 5035 1120 5957 1121
rect 5035 200 5036 1120
rect 5956 200 5957 1120
rect 5035 199 5957 200
rect 4612 -148 4716 148
rect 3423 -200 4345 -199
rect 3423 -1120 3424 -200
rect 4344 -1120 4345 -200
rect 3423 -1121 4345 -1120
rect 3000 -1320 3104 -1172
rect 3832 -1320 3936 -1121
rect 4612 -1172 4632 -148
rect 4696 -1172 4716 -148
rect 5444 -199 5548 199
rect 6224 148 6244 1172
rect 6308 148 6328 1172
rect 7056 1121 7160 1320
rect 7836 1172 7940 1320
rect 6647 1120 7569 1121
rect 6647 200 6648 1120
rect 7568 200 7569 1120
rect 6647 199 7569 200
rect 6224 -148 6328 148
rect 5035 -200 5957 -199
rect 5035 -1120 5036 -200
rect 5956 -1120 5957 -200
rect 5035 -1121 5957 -1120
rect 4612 -1320 4716 -1172
rect 5444 -1320 5548 -1121
rect 6224 -1172 6244 -148
rect 6308 -1172 6328 -148
rect 7056 -199 7160 199
rect 7836 148 7856 1172
rect 7920 148 7940 1172
rect 8668 1121 8772 1320
rect 9448 1172 9552 1320
rect 8259 1120 9181 1121
rect 8259 200 8260 1120
rect 9180 200 9181 1120
rect 8259 199 9181 200
rect 7836 -148 7940 148
rect 6647 -200 7569 -199
rect 6647 -1120 6648 -200
rect 7568 -1120 7569 -200
rect 6647 -1121 7569 -1120
rect 6224 -1320 6328 -1172
rect 7056 -1320 7160 -1121
rect 7836 -1172 7856 -148
rect 7920 -1172 7940 -148
rect 8668 -199 8772 199
rect 9448 148 9468 1172
rect 9532 148 9552 1172
rect 10280 1121 10384 1320
rect 11060 1172 11164 1320
rect 9871 1120 10793 1121
rect 9871 200 9872 1120
rect 10792 200 10793 1120
rect 9871 199 10793 200
rect 9448 -148 9552 148
rect 8259 -200 9181 -199
rect 8259 -1120 8260 -200
rect 9180 -1120 9181 -200
rect 8259 -1121 9181 -1120
rect 7836 -1320 7940 -1172
rect 8668 -1320 8772 -1121
rect 9448 -1172 9468 -148
rect 9532 -1172 9552 -148
rect 10280 -199 10384 199
rect 11060 148 11080 1172
rect 11144 148 11164 1172
rect 11892 1121 11996 1320
rect 12672 1172 12776 1320
rect 11483 1120 12405 1121
rect 11483 200 11484 1120
rect 12404 200 12405 1120
rect 11483 199 12405 200
rect 11060 -148 11164 148
rect 9871 -200 10793 -199
rect 9871 -1120 9872 -200
rect 10792 -1120 10793 -200
rect 9871 -1121 10793 -1120
rect 9448 -1320 9552 -1172
rect 10280 -1320 10384 -1121
rect 11060 -1172 11080 -148
rect 11144 -1172 11164 -148
rect 11892 -199 11996 199
rect 12672 148 12692 1172
rect 12756 148 12776 1172
rect 12672 -148 12776 148
rect 11483 -200 12405 -199
rect 11483 -1120 11484 -200
rect 12404 -1120 12405 -200
rect 11483 -1121 12405 -1120
rect 11060 -1320 11164 -1172
rect 11892 -1320 11996 -1121
rect 12672 -1172 12692 -148
rect 12756 -1172 12776 -148
rect 12672 -1320 12776 -1172
<< properties >>
string FIXED_BBOX 11404 120 12484 1200
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5.0 l 5.0 val 53.8 carea 2.00 cperi 0.19 nx 16 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1754942115
<< metal3 >>
rect -686 1172 686 1200
rect -686 148 602 1172
rect 666 148 686 1172
rect -686 120 686 148
rect -686 -148 686 -120
rect -686 -1172 602 -148
rect 666 -1172 686 -148
rect -686 -1200 686 -1172
<< via3 >>
rect 602 148 666 1172
rect 602 -1172 666 -148
<< mimcap >>
rect -646 1120 354 1160
rect -646 200 -606 1120
rect 314 200 354 1120
rect -646 160 354 200
rect -646 -200 354 -160
rect -646 -1120 -606 -200
rect 314 -1120 354 -200
rect -646 -1160 354 -1120
<< mimcapcontact >>
rect -606 200 314 1120
rect -606 -1120 314 -200
<< metal4 >>
rect -198 1121 -94 1320
rect 582 1172 686 1320
rect -607 1120 315 1121
rect -607 200 -606 1120
rect 314 200 315 1120
rect -607 199 315 200
rect -198 -199 -94 199
rect 582 148 602 1172
rect 666 148 686 1172
rect 582 -148 686 148
rect -607 -200 315 -199
rect -607 -1120 -606 -200
rect 314 -1120 315 -200
rect -607 -1121 315 -1120
rect -198 -1320 -94 -1121
rect 582 -1172 602 -148
rect 666 -1172 686 -148
rect 582 -1320 686 -1172
<< properties >>
string FIXED_BBOX -686 120 394 1200
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5.0 l 5.0 val 53.8 carea 2.00 cperi 0.19 nx 1 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
